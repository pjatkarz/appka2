���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK
��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak�et�b�n_features_in_�K
�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h2�f8�����R�(KhNNNNJ����J����K t�b�C              �?�t�bhRh&�scalar���hMC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���K
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hK�
node_count�K��nodes�h(h+K ��h-��R�(KK���h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h~hMK ��hhMK��h�hMK��h�h^K��h�h^K ��h�hMK(��h�h^K0��uK8KKt�b�Bx6         ~       	          ����?j8je3�?�           ��@       !                    _@dP,k|��?�            �v@                           �?�H�a��?8            @U@                           �?D^��#��?            �D@                          �]@f���M�?             ?@                          �f@����X�?             @������������������������       �                      @������������������������       �                     @	                          �l@      �?             8@
                          �k@      �?             0@                           �E@�θ�?             *@������������������������       �                     �?                            J@r�q��?
             (@������������������������       �                     @                           �L@����X�?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @                           @G@z�G�z�?             $@������������������������       �                      @������������������������       �                      @                          �k@�Ra����?             F@������������������������       �                     A@                           �?      �?	             $@������������������������       �                      @                           @\@      �?              @                          �n@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @"       #       	          ���ٿTc� �?�            �q@������������������������       �                     @$       c                   pq@�	�3�	�?�            @q@%       ,                   @E@ڢPRM�?�            `j@&       +                    �?�n_Y�K�?	             *@'       *                    �?����X�?             @(       )                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @-       <                   `]@ ���3�?|            �h@.       5                    �?�q�q�?             >@/       4                    o@և���X�?
             ,@0       1                    �?���!pc�?             &@������������������������       �                     @2       3                   Pb@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @6       ;                    \@      �?
             0@7       :                   �a@��S�ۿ?	             .@8       9                   @m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?=       ^                    �?�����?h             e@>       O                    �?��S�ۿ?`            �b@?       N                   �b@�T|n�q�?            �E@@       E                   �_@؇���X�?             E@A       D                   �d@�q�q�?             (@B       C                    �K@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @F       K                   �a@��S�ۿ?             >@G       H                    �? 7���B�?             ;@������������������������       �                     4@I       J                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?L       M                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?P       [                    @ 5x ��?E            �Z@Q       Z                   �l@p� V�?B            �Y@R       U                    �?h㱪��?%            �K@S       T                   �c@؇���X�?             @������������������������       �                     �?������������������������       �                     @V       Y                   �a@@��8��?!             H@W       X                    �L@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?������������������������       �                     =@������������������������       �                     H@\       ]                   �d@      �?             @������������������������       �                     @������������������������       �                     �?_       b                   0a@�q�q�?             2@`       a                   `a@      �?             (@������������������������       �                     @������������������������       �                     @������������������������       �                     @d       s                    �?�G\�c�?)            @P@e       r                    �?��X��?             <@f       k                   �_@��H�}�?             9@g       h                    �H@�8��8��?             (@������������������������       �                      @i       j                   �^@      �?             @������������������������       �                     �?������������������������       �                     @l       q                   8|@�n_Y�K�?             *@m       n                   �a@���!pc�?             &@������������������������       �                     @o       p                   �v@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @t       }                   �d@���@��?            �B@u       |                   �c@b�h�d.�?            �A@v       {                    �?      �?             0@w       x                   �`@�q�q�?             .@������������������������       �                     @y       z                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@������������������������       �                      @       �                   �b@
,UP��?�             w@�       �                    @8EGr��?�            �r@�       �                   {@�0����?�            �q@�       �                    �?4_�����?�            �q@�       �                    �R@@�s��?�            @l@�       �                   `_@�8��!�?�             l@�       �       	          ����?��7�K¨?S            @^@�       �                    �?�8��8��?             B@������������������������       �                      @�       �                   �X@г�wY;�?             A@�       �                   �g@�C��2(�?             &@������������������������       �                      @�       �                   @^@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@������������������������       �        ;            @U@�       �                   �[@,�T�6�?=             Z@�       �                    �D@8����?             7@������������������������       �                     @�       �                   0b@j���� �?	             1@�       �       	             �?�q�q�?             .@�       �                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �a@ףp=
�?             $@������������������������       �                      @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @M@H�!b	�?1            @T@�       �                   ``@ qP��B�?            �E@�       �                   Pl@��S�ۿ?             .@������������������������       �                     &@�       �       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@�       �                    @N@�˹�m��?             C@�       �                   P`@z�G�z�?             $@������������������������       �                     @�       �                    �?�q�q�?             @�       �       	          ���@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �l@h�����?             <@�       �       	          033@ףp=
�?             $@������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             2@������������������������       �                     �?�       �       	             �?�k�'7��?!            �L@������������������������       �                     �?�       �                    �?�X�C�?              L@�       �                    �?�X����?             6@�       �                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          `ff�?�d�����?             3@�       �                    [@      �?             $@������������������������       �                     @�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@�       �                   �`@�IєX�?             A@������������������������       �                     :@�       �                    �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?և���X�?             ,@������������������������       �                     @�       �                    �?z�G�z�?             $@������������������������       �                     �?�       �                   @_@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       	             @      �?+             Q@�       �                    �?��H�}�?              I@�       �                    �M@z�G�z�?             .@�       �                    �?և���X�?             @������������������������       �                     �?�       �                   �`@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �       	          ����?b�h�d.�?            �A@�       �       	          `ff�?�q�q�?             "@�       �                   �d@z�G�z�?             @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �d@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @K@ȵHPS!�?             :@������������������������       �        
             0@�       �                   �L@�z�G��?             $@������������������������       �                      @�       �                    �L@      �?              @������������������������       �                     @�       �                   @`@      �?             @�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   g@�����H�?             2@�       �                    @O@�IєX�?
             1@������������������������       �                     *@�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�t�b�values�h(h+K ��h-��R�(KK�KK��h^�B�       Ps@     �z@     @n@      _@      ;@      M@      6@      3@      4@      &@       @      @       @                      @      2@      @      $@      @      $@      @              �?      $@       @      @              @       @      �?       @               @      �?              @                      @       @               @       @       @                       @      @     �C@              A@      @      @       @              @      @      @       @      @                       @              @     �j@     �P@              @     �j@     �N@      f@      A@      @       @      @       @      @      �?              �?      @                      �?              @     �e@      :@      4@      $@      @       @      @       @              @      @      @      @                      @      @              ,@       @      ,@      �?      �?      �?      �?                      �?      *@                      �?      c@      0@     �a@      $@      B@      @      B@      @       @      @      @      @              @      @              @              <@       @      :@      �?      4@              @      �?      @                      �?       @      �?              �?       @                      �?      Z@      @     @Y@       @     �J@       @      @      �?              �?      @             �G@      �?      2@      �?      2@                      �?      =@              H@              @      �?      @                      �?      (@      @      @      @      @                      @      @              C@      ;@      "@      3@      "@      0@      �?      &@               @      �?      @      �?                      @       @      @       @      @      @              �?      @              @      �?                       @              @      =@       @      =@      @      $@      @      $@      @      @              @      @      @                      @              �?      3@                       @     �P@     �r@     �@@     �p@      ;@     0p@      9@      p@      .@     `j@      ,@     `j@      @     �]@      @     �@@       @              �?     �@@      �?      $@               @      �?       @              �?      �?      �?              �?      �?                      7@             @U@      &@     @W@      @      0@              @      @      $@      @      $@      @      �?      @                      �?      �?      "@               @      �?      �?      �?                      �?       @              @     @S@      �?      E@      �?      ,@              &@      �?      @      �?                      @              <@      @     �A@       @       @              @       @      @      �?      @      �?                      @      �?              �?      ;@      �?      "@              @      �?      @              @      �?                      2@      �?              $@     �G@      �?              "@     �G@      @      .@       @      �?              �?       @              @      ,@      @      @              @      @       @      @                       @              "@       @      @@              :@       @      @              @       @               @      �?       @                      �?      @       @      @               @       @      �?              �?       @      �?                       @      A@      A@      @@      2@      @      (@      @      @      �?               @      @              @       @                       @      =@      @      @      @      @      �?      �?      �?      �?                      �?      @               @       @       @                       @      7@      @      0@              @      @               @      @      �?      @              @      �?      �?      �?      �?                      �?       @               @      0@      �?      0@              *@      �?      @              @      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B9         x       	          ����?4�5����?�           ��@       7                   �`@�N2��?�            �w@                          �e@8�A�0��?H            �[@                           `@���N8�?             E@                           �?�S����?             C@                          �T@�+e�X�?             9@                           `R@      �?             8@       	                    �D@؇���X�?             5@������������������������       �                     �?
                          �Z@ףp=
�?             4@������������������������       �                      @                          @_@r�q��?	             (@������������������������       �                     @                           �?      �?              @������������������������       �                     �?                           `@����X�?             @������������������������       �                     �?                           @N@r�q��?             @                          @^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     @       (                    �?�������?-             Q@                           �?�X���?             F@������������������������       �                     "@       %                    �?և���X�?            �A@                            �?�㙢�c�?             7@������������������������       �                      @!       $                    �G@�����?             5@"       #                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             0@&       '                    @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?)       ,                   (p@      �?             8@*       +       	          hff�?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?-       2                    �?�q�q�?             (@.       1                   q@r�q��?             @/       0                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @3       6                   Pu@�q�q�?             @4       5                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?8       =                   @E@V��T���?�            �p@9       <                    \@@4և���?
             ,@:       ;                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@>       U                    �?������?�            �o@?       B                    �?X���[�?(            �R@@       A                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?C       H                    �?N1���?"            �N@D       G                   �`@�E��ӭ�?	             2@E       F                   �f@     ��?             0@������������������������       �                     *@������������������������       �                     @������������������������       �                      @I       J                    @D@8�$�>�?            �E@������������������������       �                      @K       P                   ``@z�G�z�?            �A@L       M                    g@�z�G��?             4@������������������������       �                     @N       O                    �?և���X�?             ,@������������������������       �                      @������������������������       �                     @Q       R                     M@��S�ۿ?
             .@������������������������       �                     (@S       T                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?V       w                   @g@L�'��T�?i            @f@W       l                    @L@ >�֕�?h            �e@X       a                    �? ��֛�?W            @b@Y       `                   �a@����ȫ�?2            �T@Z       _                    �?�����H�?             "@[       \                   Pa@؇���X�?             @������������������������       �                     @]       ^                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        +            @R@b       k                   `]@      �?%             P@c       j                   `\@z�G�z�?             $@d       i                   @[@�����H�?             "@e       f                    �F@z�G�z�?             @������������������������       �                     @g       h                   @Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     K@m       n                    �?>���Rp�?             =@������������������������       �                     $@o       r                   Hp@p�ݯ��?             3@p       q                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?s       v                   �q@؇���X�?             @t       u                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @y       �                    �?61���r�?�            Pv@z       �                    �?N1���?&            �N@{       �                    �?����X�?            �A@|       }                   �Z@�n_Y�K�?             :@������������������������       �                     @~       �                   �m@\X��t�?             7@       �                   �e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   `\@�q�q�?
             2@������������������������       �                      @�       �                   �q@      �?	             0@������������������������       �                     @�       �                    �?���Q��?             $@�       �                    b@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?�       �       	          ���@�q�q�?             @�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �H@ȵHPS!�?             :@�       �                    �?�q�q�?             @������������������������       �                      @�       �       	          033�?      �?             @������������������������       �                      @������������������������       �                      @�       �                    \@P���Q�?             4@�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@�       �                    @E@P�0�e��?�            �r@�       �                    �?���Q��?             4@�       �                    �?�8��8��?             (@������������������������       �                     "@�       �                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �l@      �?              @������������������������       �                     @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�                         pv@�	��X�?�            @q@�       �                   P`@�t�o}�?�            q@�       �       	          `ff@     ��?M             `@�       �                   Ph@����?E            @\@�       �       	          033�?�}�+r��?             C@������������������������       �                     2@�       �                    �?ףp=
�?             4@�       �                    W@؇���X�?	             ,@������������������������       �                     �?�       �                    �?$�q-�?             *@�       �       	              @؇���X�?             @�       �                   `_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?��n�?+            �R@�       �                   �[@H%u��?             9@�       �                   `n@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �j@�}�+r��?             3@�       �       	          pff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             0@�       �                    �?H.�!���?             I@�       �                    �?������?            �B@������������������������       �                     @�       �                   0i@�r����?             >@������������������������       �                      @�       �                   �`@@4և���?             <@������������������������       �                     6@�       �                    �?�q�q�?             @������������������������       �                     @�       �                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �[@��
ц��?             *@������������������������       �                      @�       �                   �\@���|���?             &@������������������������       �                      @�       �                   �b@�<ݚ�?             "@�       �       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	             
@�q�q�?             .@�       �                    �?�n_Y�K�?             *@�       �                    �?�����H�?             "@�       �                   8p@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�������?b             b@�       �                   `b@�t����?             1@������������������������       �                     (@�       �                   �d@���Q��?             @�       �                   `o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�                          �R@     ��?U             `@�       �       	          ����?��b�h8�?T            �_@�       �                    �?z�G�z�?             9@�       �                    �K@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?      �?             0@�       �                   ``@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     @�                          �c@г�wY;�?F            �Y@�       �       	          ����?p���?D             Y@�       �                   �Q@������?            �D@�       �                     N@r�q��?             (@�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     =@������������������������       �        *            �M@                        �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h^�BP       �t@     y@     p@      ^@     �F@     @P@      $@      @@      @      @@      @      3@      @      2@      @      2@      �?               @      2@               @       @      $@              @       @      @              �?       @      @      �?              �?      @      �?       @      �?                       @              @      @                      �?              *@      @             �A@     �@@      =@      .@      "@              4@      .@      3@      @               @      3@       @      @       @               @      @              0@              �?      &@              &@      �?              @      2@      �?      &@              &@      �?              @      @      �?      @      �?       @               @      �?                      @      @       @      @      �?      @                      �?              �?     �j@     �K@      �?      *@      �?       @      �?                       @              &@     `j@      E@      G@      =@      *@      �?      *@                      �?     �@@      <@      @      *@      @      *@              *@      @               @              <@      .@               @      <@      @      ,@      @      @               @      @       @                      @      ,@      �?      (@               @      �?       @                      �?     �d@      *@     �d@      $@     �a@      @     @T@      �?       @      �?      @      �?      @               @      �?              �?       @               @             @R@              O@       @       @       @       @      �?      @      �?      @              �?      �?      �?                      �?      @                      �?      K@              6@      @      $@              (@      @      &@      �?      &@                      �?      �?      @      �?       @               @      �?                      @              @      S@     �q@     �@@      <@      $@      9@      $@      0@              @      $@      *@      @      �?              �?      @              @      (@       @              @      (@              @      @      @      @      @      @                      @      �?      @              �?      �?       @      �?      �?              �?      �?                      �?              "@      7@      @      @       @       @               @       @               @       @              3@      �?      �?      �?              �?      �?              2@             �E@     �o@       @      (@      �?      &@              "@      �?       @      �?                       @      @      �?      @              @      �?      @                      �?     �A@      n@      @@      n@      5@     �Z@      0@     @X@       @      B@              2@       @      2@       @      (@      �?              �?      (@      �?      @      �?      @              @      �?                       @              @              @      ,@     �N@      @      6@       @      @       @                      @      �?      2@      �?       @      �?                       @              0@      &@     �C@      @     �@@              @      @      :@       @               @      :@              6@       @      @              @       @      �?       @                      �?      @      @               @      @      @               @      @       @      @       @      @                       @      @              @      $@      @       @      �?       @      �?      @               @      �?      �?              �?      �?                      @      @                       @      &@     �`@       @      .@              (@       @      @       @      �?       @                      �?               @      "@     �]@       @     �]@      @      4@      @      @      @                      @       @      ,@       @      &@              &@       @                      @      @     �X@       @     �X@       @     �C@       @      $@       @       @       @                       @               @              =@             �M@      �?      �?      �?                      �?      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK녔h}�Bh3         2                    �?p�Vv���?�           ��@              	          ����?�>�p���?Y             b@                          �Q@�����H�?4            @T@                          a@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?�:�^���?1            �S@                           d@�t����?
             1@	       
                     J@8�Z$���?             *@������������������������       �                      @                           ]@���Q��?             @������������������������       �                      @                           �?�q�q�?             @                          �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                          @d@      �?             @������������������������       �                     @������������������������       �                     �?                           �?�]0��<�?'            �N@������������������������       �        "             J@                           �L@�<ݚ�?             "@                           a@�q�q�?             @                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       -                    �?     ��?%             P@       $                    �?������?            �F@        !                   �R@j���� �?             1@������������������������       �                     @"       #       	          `ff@����X�?             ,@������������������������       �                     $@������������������������       �                     @%       ,       	          ����?@4և���?             <@&       '                    �?"pc�
�?             &@������������������������       �                     @(       )                   �m@����X�?             @������������������������       �                     �?*       +                   @_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@.       1       	          ����?�}�+r��?             3@/       0                   `c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@3       �                    �?~�.���?�           h�@4       ?                   �_@|�38���?�            �t@5       6                    �?���J��?C            �Y@������������������������       �        -            @Q@7       8       	          033�?�FVQ&�?            �@@������������������������       �                     9@9       :                   @`@      �?              @������������������������       �                     �?;       >                    �?؇���X�?             @<       =                   `]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@       s                    �?P̏����?�            �l@A       T                   �`@�i#[��?9             U@B       O                   �k@8^s]e�?             =@C       F                   �Y@���Q��?             4@D       E                    �?����X�?             @������������������������       �                     @������������������������       �                      @G       L                    �?�θ�?
             *@H       K                   pi@ףp=
�?             $@I       J                   �g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @M       N                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?P       S                    �G@�����H�?             "@Q       R                   Hy@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @U       l                   �n@N{�T6�?#            �K@V       g                   �e@���y4F�?             C@W       Z                    �D@6YE�t�?            �@@X       Y       	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @[       f                   pk@ףp=
�?             >@\       e       	          hff�?r�q��?
             2@]       d                    �?�t����?	             1@^       c       	          ����?�r����?             .@_       `                   �b@"pc�
�?             &@������������������������       �                     @a       b                   �\@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@h       i                    �D@���Q��?             @������������������������       �                      @j       k                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @m       r                   b@������?             1@n       q                   �z@�q�q�?             @o       p                    @N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@t       �                   (q@�5?,R�?b             b@u       �                   q@0w-!��?F             Y@v       �                    �?�^'�ë�?E            @X@w       �                   �e@      �?6             T@x       y                   i@���!���?5            �S@������������������������       �                     2@z       �                   @j@f>�cQ�?(            �N@{       |       	             �?����X�?             @������������������������       �                     �?}       �                   �i@r�q��?             @~              	          033�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �       	            �?�>����?#             K@�       �       	          ����?      �?             @�       �                   `a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �[@`2U0*��?              I@������������������������       �                     ,@�       �                    �J@�X�<ݺ?             B@�       �                    @J@�r����?             .@�       �                   �m@$�q-�?	             *@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@������������������������       �                     �?������������������������       �                     1@������������������������       �                     @������������������������       �                     F@�       �       	          ����?��?�            0p@�       �                    @�}���?x             h@�       �                   �X@,�"���?l            @e@�       �                    @G@���!pc�?	             &@������������������������       �                      @�       �                   @`@�����H�?             "@�       �                   `V@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �O@���C��?c            �c@�       �                    �?      �?              @������������������������       �                      @�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �K@tX�}}��?]            �b@�       �                   �g@���#�İ?F            �]@�       �                    @H@ ���J��?E            @]@�       �                    �G@xL��N�?+            �R@�       �                   �a@����e��?&            �P@�       �                   `a@��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                    �I@�       �                   �d@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                    �E@������������������������       �                     �?�       �                   �a@�q�q�?            �@@�       �       	          ����?�G�z��?             4@�       �                    �?�q�q�?             .@�       �                   �i@X�<ݚ�?             "@������������������������       �                      @�       �                   �a@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    @L@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@�       �                   �c@�û��|�?             7@�       �                   �p@��.k���?	             1@�       �                   `Q@      �?             (@������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                     @�       �                   P`@r�q��?0            �P@�       �                    `@�LQ�1	�?             7@�       �       	          ��� @�d�����?             3@�       �                   �^@�eP*L��?
             &@�       �                   �o@����X�?             @�       �                   �\@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	             @      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     E@Du9iH��?            �E@������������������������       �                     �?�       �                   pb@���N8�?             E@������������������������       �                    �@@�       �                   �h@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       @t@     �y@     �Y@     �E@      R@      "@      �?       @      �?                       @     �Q@      @      (@      @      &@       @       @              @       @       @              �?       @      �?      �?              �?      �?                      �?      �?      @              @      �?             �M@       @      J@              @       @      @       @      @      �?      @                      �?              �?      @              >@      A@      (@     �@@      $@      @              @      $@      @      $@                      @       @      :@       @      "@              @       @      @      �?              �?      @      �?                      @              1@      2@      �?      @      �?      @                      �?      .@             �k@     �v@      M@      q@       @      Y@             @Q@       @      ?@              9@       @      @      �?              �?      @      �?      @              @      �?                      @      L@     �e@     �E@     �D@      "@      4@       @      (@      @       @      @                       @      @      $@      �?      "@      �?      �?              �?      �?                       @       @      �?       @                      �?      �?       @      �?       @      �?                       @              @      A@      5@      >@       @      <@      @      �?       @      �?                       @      ;@      @      .@      @      .@       @      *@       @      "@       @      @              @       @      @                       @      @               @                      �?      (@               @      @               @       @      �?              �?       @              @      *@      @       @      @      �?      @                      �?              �?              &@      *@     ``@      *@     �U@      $@     �U@      $@     �Q@      "@     �Q@              2@      "@      J@      @       @              �?      @      �?      @      �?      @                      �?       @              @      I@       @       @      �?       @               @      �?              �?               @      H@              ,@       @      A@       @      *@      �?      (@               @      �?      @              @      �?              �?      �?              �?      �?                      5@      �?                      1@      @                      F@     �d@     �W@      c@      D@      b@      :@      @       @       @              �?       @      �?      @      �?      �?      �?                      �?              @              @     �a@      2@      @      @       @              @      @              @      @              a@      .@     �\@      @     �\@      @     �Q@      @     @P@      �?      ,@      �?      ,@                      �?     �I@              @       @      @                       @     �E@                      �?      6@      &@      "@      &@      @      $@      @      @               @      @      @      @                      @      �?      @      �?                      @      @      �?      @                      �?      *@              "@      ,@      "@       @      "@      @              @      "@                      @              @      &@     �K@       @      .@      @      ,@      @      @       @      @       @       @              �?       @      �?      �?              �?      �?              �?      �?                      @      @      �?              �?      @                       @      @      �?       @              �?      �?              �?      �?              @      D@      �?               @      D@             �@@       @      @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK���h}�Bx6         r                   �`@U�ք�?�           ��@       C                   �`@�~6�]�?�            @u@       "                    �?�G�z��?n             d@                           �?      �?/             Q@                           �?�"U����?%            �I@                          p`@�Q����?             D@                           �?�s��:��?             C@       	       	          ����?��S�ۿ?             .@������������������������       �        	             (@
                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?8����?             7@                           [@$�q-�?             *@                          �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             &@                          �Z@���Q��?             $@������������������������       �                     @                          �Y@؇���X�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     &@                           �?�t����?
             1@������������������������       �                     �?              	          ����?      �?	             0@������������������������       �                     "@        !                    �L@؇���X�?             @������������������������       �                     @������������������������       �                     �?#       B                    `@��A��??             W@$       3                   �^@z���=��?4            @S@%       (                    [@@4և���?             E@&       '       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       0                   Hs@�7��?            �C@*       +                    @L@��?^�k�?            �A@������������������������       �                     5@,       /                    \@@4և���?
             ,@-       .                    Y@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@1       2                   �t@      �?             @������������������������       �                     �?������������������������       �                     @4       7                    �?����X�?            �A@5       6                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @8       ?       	          ����?V�a�� �?             =@9       :                   �Y@�n_Y�K�?             *@������������������������       �                     @;       <       	          ����?      �?              @������������������������       �                      @=       >                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?@       A                   @_@      �?	             0@������������������������       �                     �?������������������������       �                     .@������������������������       �                     .@D       M                    �G@4?,R��?k            �f@E       F                   @a@�z�G��?             $@������������������������       �                     �?G       H                    �?�<ݚ�?             "@������������������������       �                     @I       J                    �?      �?             @������������������������       �                     �?K       L                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @N       c       	          033�?�̨�`<�?d            @e@O       b                    �?      �?             F@P       _       	          ����?��>4և�?             <@Q       ^                     O@���!pc�?             6@R       Y                    �?���Q��?
             .@S       T                    �?�����H�?             "@������������������������       �                     @U       X                    �?r�q��?             @V       W                     K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Z       [                    �?r�q��?             @������������������������       �                     @\       ]                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @`       a                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             0@d       q                    `R@�X�<ݺ?I            �_@e       j                    `@`J����?H            �^@f       g                    @@���a��?C            �\@������������������������       �        A            �[@h       i                    �?      �?             @������������������������       �                     �?������������������������       �                     @k       p                    @N@      �?              @l       m       	          ����?      �?             @������������������������       �                      @n       o       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @s       �                    �?�����?           �x@t       �                    @L@�z�G��?�            �t@u       �       	             @���0��?�            �m@v       �                   @g@B�Y��f�?�            �l@w       �                   �`@&^�r���?�            @l@x       �                   `]@�Z��=��?j            �c@y       z                   pb@      �?             D@������������������������       �                     .@{       |                   0c@���Q��?             9@������������������������       �                     @}       �                   �p@�X����?             6@~                           �?     ��?             0@������������������������       �                     @�       �                   �i@�z�G��?             $@������������������������       �                     @�       �                    �F@      �?             @������������������������       �                      @�       �                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?|�űN�?P            @]@������������������������       �                     F@�       �                    �G@L������?5            @R@�       �                    �?���N8�?             E@������������������������       �                     �?�       �                    @��Y��]�?            �D@������������������������       �                     D@������������������������       �                     �?�       �                    �?�n`���?             ?@�       �                   �^@      �?
             (@�       �                    b@z�G�z�?             @������������������������       �                      @�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `@����X�?             @������������������������       �                     @�       �       	          433�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     3@�       �                   �`@�G�5��?1            @Q@�       �                   @c@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    @Z���c��?,            �O@�       �                    �?�:�B��?)            �M@������������������������       �                     &@�       �       	          @33�?�q�q�?"             H@�       �                   �f@�C��2(�?            �@@�       �                   xp@`Jj��?             ?@������������������������       �                     2@�       �                    �?8�Z$���?             *@�       �                   �p@�8��8��?
             (@�       �                    @E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�       �                   g@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?��S���?             .@������������������������       �                      @�       �                    �G@�n_Y�K�?             *@������������������������       �                     @�       �                     J@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �                   `f@      �?             @�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?z�G�z�?	             $@������������������������       �                     �?�       �                   n@�����H�?             "@������������������������       �                     @�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �j@��c:�?7             W@�       �                   @a@     ��?             0@������������������������       �                      @�       �                    @N@      �?              @������������������������       �                     @������������������������       �                     @�       �       	          `ff�?���=A�?+             S@�       �                    �?*O���?             B@�       �       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �q@������?             >@�       �                    �?؇���X�?             5@������������������������       �                     "@�       �                    �M@      �?             (@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?X�<ݚ�?             "@������������������������       �                     @�       �                   0b@�q�q�?             @������������������������       �                      @�       �                   ht@      �?             @������������������������       �                     �?�       �                   u@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?P���Q�?             D@������������������������       �                     >@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �?     ��?)             P@������������������������       �                     B@�       �                   �o@��X��?             <@�       �                    @z�G�z�?             4@�       �                   �O@�S����?             3@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @M@      �?             0@������������������������       �                     (@�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �q@      �?              @������������������������       �                     @�       �                   c@      �?             @������������������������       �                     �?������������������������       �                     @�t�b�l!     h�h(h+K ��h-��R�(KK�KK��h^�B�        t@     �y@      R@     �p@     �G@     @\@      A@      A@      @@      3@      5@      3@      5@      1@      ,@      �?      (@               @      �?              �?       @              @      0@      �?      (@      �?      �?      �?                      �?              &@      @      @              @      @      �?      �?      �?              �?      �?              @                       @      &@               @      .@      �?              �?      .@              "@      �?      @              @      �?              *@     �S@      *@      P@      @     �C@      �?       @      �?                       @       @     �B@      �?      A@              5@      �?      *@      �?      @              @      �?                      $@      �?      @      �?                      @      $@      9@      @       @               @      @              @      7@      @       @              @      @      @               @      @      �?      @                      �?      �?      .@      �?                      .@              .@      9@     `c@      @      @              �?      @       @      @               @       @              �?       @      �?              �?       @              2@      c@      &@     �@@      &@      1@      @      0@      @      "@      �?       @              @      �?      @      �?       @               @      �?                      @      @      �?      @               @      �?       @                      �?              @      @      �?              �?      @                      0@      @     �]@      @     �]@      �?     �\@             �[@      �?      @      �?                      @      @      @      @      �?       @              �?      �?              �?      �?                      @      @             @o@      b@     �l@     �X@      h@     �F@     �g@     �B@     �g@     �A@     `a@      2@      >@      $@      .@              .@      $@              @      .@      @      "@      @      @              @      @              @      @      @       @              �?      @      �?                      @      @             @[@       @      F@             @P@       @      D@       @              �?      D@      �?      D@                      �?      9@      @      @      @      @      �?       @               @      �?       @                      �?       @      @              @       @      �?       @                      �?      3@              J@      1@       @      @              @       @              I@      *@     �H@      $@      &@              C@      $@      >@      @      =@       @      2@              &@       @      &@      �?      �?      �?      �?                      �?      $@                      �?      �?      �?              �?      �?               @      @               @       @      @      @              @      @              @      @              �?      @      �?      �?              �?      �?                       @               @       @       @      �?              �?       @              @      �?      �?      �?                      �?      C@      K@      *@      @       @              @      @      @                      @      9@     �I@      7@      *@      �?      @              @      �?              6@       @      2@      @      "@              "@      @      �?      @              @      �?               @              @      @              @      @       @       @               @       @      �?              �?       @               @      �?               @      C@              >@       @       @       @                       @      3@     �F@              B@      3@      "@      0@      @      0@      @      �?       @               @      �?              .@      �?      (@              @      �?              �?      @                      �?      @      @              @      @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuM	hvh(h+K ��h-��R�(KM	��h}�B�9         �       	          ����?4�5����?�           ��@       7                    @J@�Ff��K�?�            x@                           �?H芦��?�            �j@                          i@J�����?/            @S@                           �?��� ��?             ?@                          �Z@��s����?             5@������������������������       �                      @       	                     H@�KM�]�?
             3@������������������������       �                     .@
                           @I@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     $@                            B@���j��?             G@������������������������       �                     @                          �Z@>��C��?            �E@������������������������       �                     @                          hp@z�G�z�?             D@                          �Y@�>����?             ;@                           l@      �?              @������������������������       �                     �?������������������������       �                     �?                          �b@`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?                          �a@�n_Y�K�?             *@������������������������       �                     @                          0d@r�q��?             @������������������������       �                     @������������������������       �                     �?                            �?���.�6�?W            @a@������������������������       �                    �G@!       .                   `]@�ɮ����?<            �V@"       -                   `\@�q�q�?
             .@#       ,                    �?����X�?	             ,@$       %       	          ������	j*D�?             *@������������������������       �                     �?&       +                   �o@�q�q�?             (@'       *                   @[@�����H�?             "@(       )                    i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?/       0                   `a@�}�+r��?2             S@������������������������       �                     F@1       2                   �b@      �?             @@������������������������       �                     &@3       4                   �d@��s����?             5@������������������������       �                     @5       6                   pe@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@8       o                    �?k�q��?s            @e@9       F                   �a@�������?S             ]@:       C                    �?8����?             7@;       @                   �_@���Q��?             .@<       =                   �`@�����H�?             "@������������������������       �                     @>       ?                    �?      �?              @������������������������       �                     �?������������������������       �                     �?A       B                    @r�q��?             @������������������������       �                     @������������������������       �                     �?D       E                   �`@      �?              @������������������������       �                     @������������������������       �                     �?G       n                   �g@��!���?D            @W@H       O                    �?@S�)�q�?C            �V@I       N                    �?�g�y��?             ?@J       K                   d@�����H�?             "@������������������������       �                     @L       M                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     6@P       m                   xt@������?/             N@Q       ^                    �?>���Rp�?.             M@R       U                   �\@\X��t�?             7@S       T                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?V       ]       	          @33�?�t����?             1@W       X                   �f@�eP*L��?	             &@������������������������       �                      @Y       Z                   @^@X�<ݚ�?             "@������������������������       �                     @[       \                   �n@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @_       d                    b@(N:!���?            �A@`       a       	          pff�?`2U0*��?             9@������������������������       �                     4@b       c                     L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?e       l                   �p@�z�G��?	             $@f       g                    X@�<ݚ�?             "@������������������������       �                     �?h       k                   c@      �?              @i       j                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @p       �                   �b@�{��?��?              K@q       v                    �?8��8���?             H@r       u                   �^@���Q��?             @s       t                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @w       |                   �`@X�EQ]N�?            �E@x       {                   �Z@ ��WV�?             :@y       z                    �O@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@}       �       	             �?������?             1@~       �                    �?؇���X�?	             ,@       �                   �T@����X�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �c@�q�q�?             @������������������������       �                      @�       �                     Q@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@�?ʵ���?�            �u@�       �       	          ����?؇���X�?�            �q@�       �                   �`@~X�<��?2             R@�       �                    �E@Z�K�D��?            �G@������������������������       �                      @�       �                    W@��Zy�?            �C@�       �                    `@�����H�?             "@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          `ff�?��S���?             >@������������������������       �                     �?�       �                   @Z@П[;U��?             =@������������������������       �                     @�       �                    �K@��H�}�?             9@�       �                   �`@և���X�?
             ,@�       �                    �?z�G�z�?             $@������������������������       �                     �?�       �                    �?�����H�?             "@�       �                   @_@r�q��?             @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                     P@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?HP�s��?             9@������������������������       �                     4@�       �                    @L@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?ܾ�z�<�?�             j@�       �                   ``@���`uӽ?k             d@�       �                    �?�y��*�?*             M@�       �                    �?���!pc�?             &@�       �                   �`@���Q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	             @dP-���?#            �G@�       �                    �?P���Q�?             D@�       �                   `_@�8��8��?             8@������������������������       �                     .@�       �                   j@�<ݚ�?             "@�       �       	             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@�       �                   �Z@����X�?             @������������������������       �                     �?�       �                   �_@r�q��?             @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   P`@ f^8���?A            �Y@�       �                   �r@����ȫ�?1            �T@������������������������       �        '            �O@�       �                    �?�}�+r��?
             3@������������������������       �        	             2@������������������������       �                     �?�       �                   p`@�����?             5@������������������������       �                     �?�       �                   �c@P���Q�?             4@������������������������       �                     0@�       �                    @O@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��|�5��?            �G@�       �                   �n@؇���X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   0g@      �?             D@�       �                    @�d�����?             3@�       �                    ]@8�Z$���?	             *@�       �                    �?�q�q�?             @������������������������       �                      @�       �                     O@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   @_@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     5@�             	             @ꮃG��?/            @Q@�       �                    �?N{�T6�?%            �K@�       �                   �g@���"͏�?            �B@������������������������       �                      @�       �                    �?z�G�z�?            �A@������������������������       �                     (@�       �                    �L@8����?             7@�       �                   �q@r�q��?             2@�       �                   �\@���!pc�?	             &@������������������������       �                      @�       �                   �e@�����H�?             "@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   pc@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�                          �?�q�q�?             2@�                           q@$�q-�?	             *@������������������������       �                     &@                        pd@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         �?@4և���?
             ,@������������������������       �                     &@                        �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM	KK��h^�B�       �t@     y@      p@     �_@     �d@     �H@     �B@      D@      @      ;@      @      1@       @               @      1@              .@       @       @       @                       @              $@     �@@      *@              @     �@@      $@              @     �@@      @      9@       @      �?      �?              �?      �?              8@      �?      8@                      �?       @      @      @              �?      @              @      �?              `@      "@     �G@             �T@      "@      $@      @      $@      @      "@      @      �?               @      @       @      �?      �?      �?      �?                      �?      @                      @      �?                      �?      R@      @      F@              <@      @      &@              1@      @              @      1@      �?              �?      1@              W@     �S@     @T@     �A@      @      0@      @      "@      �?       @              @      �?      �?              �?      �?              @      �?      @                      �?      �?      @              @      �?             �R@      3@     �R@      1@      >@      �?       @      �?      @               @      �?       @                      �?      6@              F@      0@      F@      ,@      *@      $@      �?      @              @      �?              (@      @      @      @       @              @      @      @              �?      @              @      �?              @              ?@      @      8@      �?      4@              @      �?      @                      �?      @      @      @       @              �?      @      �?      �?      �?      �?                      �?      @                      �?               @               @      &@     �E@      @     �D@       @      @       @      �?       @                      �?               @      @      C@      �?      9@      �?      @              @      �?                      2@      @      *@       @      (@       @      @       @      �?              �?       @                      @              @       @      �?       @                      �?      @       @       @               @       @       @                       @     �R@      q@      D@      n@      3@     �J@      1@      >@               @      1@      6@      �?       @              @      �?       @               @      �?              0@      ,@              �?      0@      *@              @      0@      "@      @       @       @       @      �?              �?       @      �?      @      �?      �?              �?      �?                      @              @      @              $@      �?      $@                      �?       @      7@              4@       @      @       @                      @      5@     `g@      $@     �b@      @     �I@      @       @      @       @      �?       @      �?                       @       @                      @      @     �E@       @      C@       @      6@              .@       @      @       @      �?       @                      �?              @              0@       @      @      �?              �?      @      �?      �?              �?      �?                      @      @      Y@      �?     @T@             �O@      �?      2@              2@      �?               @      3@      �?              �?      3@              0@      �?      @              @      �?              &@      B@      @      �?      @               @      �?       @                      �?      @     �A@      @      ,@       @      &@       @      @               @       @       @               @       @                      @      @      @      @                      @              5@     �A@      A@      A@      5@      <@      "@               @      <@      @      (@              0@      @      .@      @       @      @               @       @      �?      @              �?      �?      �?                      �?      @              �?      @      �?                      @      @      (@      �?      (@              &@      �?      �?      �?                      �?      @              �?      *@              &@      �?       @      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B88         �       	          ����?6������?�           ��@                          @E@��_���?�             w@       
                    �?�S����?$            �L@                           �? >�֕�?            �A@������������������������       �                     9@                           [@z�G�z�?             $@������������������������       �                     @       	                   �]@���Q��?             @������������������������       �                      @������������������������       �                     @                          �_@�X����?             6@                          `]@@4և���?             ,@������������������������       �                     "@                           �?z�G�z�?             @������������������������       �                     @                          �^@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?              @������������������������       �                     @������������������������       �                      @       W                   �n@�W�o���?�            ps@       >                    �?\[j��?v             g@       =                    �?��0u���?&             N@       $                   �]@�BbΊ�?$             M@       #                   j@      �?             0@       "                    �?z�G�z�?             $@                           @G@����X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?        !                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @%       :                   �e@r�q��?             E@&       /                   pf@�ݜ�?            �C@'       .                    �?և���X�?             @(       )                    �L@z�G�z�?             @������������������������       �                      @*       -                     O@�q�q�?             @+       ,                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @0       5                   �i@      �?             @@1       4       	          @33�?؇���X�?             @2       3                    �L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @6       7                    @O@`2U0*��?             9@������������������������       �        	             4@8       9                    �O@z�G�z�?             @������������������������       �                     �?������������������������       �                     @;       <                     F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @?       B                   �W@0{�v��?P            @_@@       A                    �?      �?             @������������������������       �                     @������������������������       �                     @C       T                    `P@hx<?v��?N            �]@D       M                   �l@ T���v�?K            @\@E       L                   �a@�q�q�??             X@F       K                   p`@Pa�	�?            �@@G       H                    �?@4և���?             ,@������������������������       �        	             (@I       J                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@������������������������       �        )            �O@N       O                    �?�t����?             1@������������������������       �                     &@P       Q                   �l@�q�q�?             @������������������������       �                     �?R       S                    @G@z�G�z�?             @������������������������       �                     @������������������������       �                     �?U       V                    �?      �?             @������������������������       �                     @������������������������       �                     @X       u                    �?X�Cc�?Q            �_@Y       Z                   �Z@�d�����?             C@������������������������       �                     �?[       b                    @F@���"͏�?            �B@\       a                    �D@�C��2(�?             &@]       `                    �?z�G�z�?             @^       _                    _@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       j                    �?�	j*D�?             :@d       e                     J@���Q��?             $@������������������������       �                     @f       g                   �b@և���X�?             @������������������������       �                      @h       i                    �?���Q��?             @������������������������       �                      @������������������������       �                     @k       n                   Xp@      �?	             0@l       m                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?o       t                   b@@4և���?             ,@p       s                    @J@z�G�z�?             @q       r                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@v       w                    Z@
�GN��?:             V@������������������������       �                     @x       �                    �K@P�;�&��?8            @U@y       ~                   `]@     ��?(             P@z       {                   �e@���|���?             &@������������������������       �                     @|       }                   p@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       �                    @�&=�w��?#            �J@�       �                    �? pƵHP�?"             J@������������������������       �                     E@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                    @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �b@�ՙ/�?             5@�       �                   ht@     ��?             0@�       �                   �`@؇���X�?             ,@�       �                    �L@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                   u@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?xƅd�?�            �v@�       �                    �? �&�T�?�            @q@�       �       	          033�?���Q��?              I@�       �                   @[@      �?             @@������������������������       �                     @�       �                    �?д>��C�?             =@�       �                   �`@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        	             4@�       �                    �?�q�q�?             2@������������������������       �                     (@������������������������       �                     @�       �                   �e@��ti�?�            @l@�       �                   P`@r�q��?�             k@�       �       	             �?�t`�4 �?J            �^@������������������������       �                     �?�       �                    @8@W"�h�?I            @^@�       �                    �?��(\���?H             ^@�       �                   �W@������?	             .@������������������������       �                     @������������������������       �                     &@�       �                   i@���N8�??            @Z@������������������������       �                    �G@�       �                    �?��ϭ�*�?&             M@�       �                    �L@4��?�?#             J@�       �                   �_@؇���X�?            �A@�       �                   pp@�q�q�?             .@�       �                    �?����X�?             @������������������������       �                     �?�       �                   @]@r�q��?             @������������������������       �                     @�       �                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     4@������������������������       �                     1@������������������������       �                     @������������������������       �                     �?�       �                    �?V��N��?<            �W@�       �                   �Z@F�t�K��?#            �L@�       �                   0a@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	          033@f1r��g�?             �J@�       �       	          033@x�����?            �C@�       �                   p`@�MI8d�?            �B@������������������������       �                     �?�       �                   pb@4?,R��?             B@�       �                    �N@�t����?             A@�       �                     M@"pc�
�?             6@�       �       	          ����?      �?
             0@�       �                   �j@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   @d@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     (@�       �                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        	             ,@�       �                   b@؀�:M�?            �B@�       �                    �H@r�q��?             @�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	             @¦	^_�?             ?@�       �                    X@�\��N��?             3@������������������������       �                      @�       �                    �L@��.k���?             1@�       �       	          ����?�<ݚ�?             "@�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@�       �                   �X@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �M@,sI�v�?6            �V@�       �       	          ����?      �?             D@������������������������       �                     @�       �                    @J@�t����?             A@������������������������       �                     .@�       �       	          ����?�\��N��?             3@�       �                    @M@�<ݚ�?             "@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?�z�G��?	             $@�       �                    e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�              	          ����?p���?             I@�       �                   �m@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �E@�t�bh�h(h+K ��h-��R�(KMKK��h^�B       �t@     �x@      o@     �]@      "@      H@       @     �@@              9@       @       @              @       @      @       @                      @      @      .@      �?      *@              "@      �?      @              @      �?      �?      �?                      �?      @       @      @                       @      n@     �Q@     �c@      :@     �E@      1@     �E@      .@       @       @       @       @       @      @              @       @      �?      �?              �?      �?              �?      �?                      @      @             �A@      @      A@      @      @      @      @      �?       @               @      �?      �?      �?              �?      �?              �?                       @      >@       @      @      �?      @      �?      @                      �?       @              8@      �?      4@              @      �?              �?      @              �?       @               @      �?                       @      ]@      "@      @      @      @                      @     @\@      @     �[@      @     �W@      �?      @@      �?      *@      �?      (@              �?      �?      �?                      �?      3@             �O@              .@       @      &@              @       @              �?      @      �?      @                      �?      @      @      @                      @     @T@     �F@      $@      <@      �?              "@      <@      �?      $@      �?      @      �?      @              @      �?                      �?              @       @      2@      @      @      @              @      @               @      @       @               @      @               @      ,@      �?      �?      �?                      �?      �?      *@      �?      @      �?       @               @      �?                       @              "@     �Q@      1@              @     �Q@      ,@      M@      @      @      @      @              �?      @      �?                      @     �I@       @     �I@      �?      E@              "@      �?      @               @      �?              �?       @                      �?      *@       @      *@      @      (@       @      @       @               @      @              "@              �?      �?              �?      �?                      @     �U@     �q@     �R@      i@      >@      4@      8@       @              @      8@      @      @      @      @                      @      4@              @      (@              (@      @             �F@     �f@      B@     �f@      &@     �[@      �?              $@     �[@      "@     �[@      @      &@      @                      &@      @      Y@             �G@      @     �J@      @     �G@      @      >@      @      $@      @       @              �?      @      �?      @               @      �?              �?       @                       @              4@              1@              @      �?              9@     @Q@      &@      G@      @      �?              �?      @               @     �F@       @      ?@      @      ?@      �?              @      ?@      @      >@      @      2@      �?      .@      �?      @              @      �?                      $@      @      @      @                      @              (@      �?      �?      �?                      �?       @                      ,@      ,@      7@      @      �?      �?      �?              �?      �?              @              "@      6@      "@      $@               @      "@       @      @       @      �?       @               @      �?              @               @      @              @       @      @       @                      @              (@      "@      �?              �?      "@              &@     �S@      $@      >@              @      $@      8@              .@      $@      "@      @       @      @      �?      @                      �?              �?      @      @      @      �?      @                      �?              @      �?     �H@      �?      @              @      �?                     �E@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK녔h}�Bh3         P                   P`@U�ք�?�           ��@       /                    �?j=M>�:�?�            �s@                           �?X�Emq�?A            �Z@                           `@r֛w���?             ?@������������������������       �                     "@                           �?���|���?
             6@������������������������       �                     @       	       	          ����?      �?             0@������������������������       �                     (@
                            P@      �?             @������������������������       �                      @������������������������       �                      @                          �\@�sly47�?/            �R@                          @X@8�Z$���?            �C@������������������������       �                     $@                           �E@V�a�� �?             =@������������������������       �                     @              	          ����?ȵHPS!�?             :@                          �Y@r�q��?             2@                           ]@      �?             @������������������������       �                      @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                      @       (                   `n@)O���?             B@       #       	          `ff�?��H�}�?             9@       "                    �H@���y4F�?             3@       !                    �?X�<ݚ�?             "@                            �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     $@$       '                    �?r�q��?             @%       &                    \@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @)       .                    �?�C��2(�?             &@*       -       	             �?�q�q�?             @+       ,                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @0       C                   P`@���ȑ��?             j@1       B                    �?ȵHPS!�?2            �S@2       5                    �?��ɉ�?*            @P@3       4       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?6       =                   `_@�8��8��?'             N@7       8                   (p@ ��WV�?!             J@������������������������       �                    �D@9       :                    @L@"pc�
�?             &@������������������������       �                      @;       <                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @>       ?                    �K@      �?              @������������������������       �                     @@       A                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@D       O                    �R@�z�N��?M            ``@E       F                   0q@ ����?L            @`@������������������������       �        <             Y@G       J                    �G@��S�ۿ?             >@H       I       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?K       N       	             �?h�����?             <@L       M                   �b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@������������������������       �                     �?Q       �       	          ��� @@<QR���?           0z@R       �                    �?*2��`B�?�            Px@S       `                    �D@6�Nӆ�?a            �b@T       _                   �r@�LQ�1	�?             7@U       ^                   �f@�C��2(�?             6@V       W                   `]@���N8�?             5@������������������������       �                     &@X       ]                   �l@ףp=
�?             $@Y       Z                   �[@      �?             @������������������������       �                      @[       \                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?a       ~                    �?P�B�y��?P            @_@b       y                   �a@�LQ�1	�?+            @Q@c       v                   ``@�BbΊ�?&             M@d       e                   `T@#z�i��?            �D@������������������������       �                     @f       m                    �?      �?             B@g       h                    �?���Q��?             .@������������������������       �                     @i       j                   `\@���Q��?             $@������������������������       �                     @k       l                   @f@�q�q�?             @������������������������       �                      @������������������������       �                     @n       u                   �s@؇���X�?             5@o       t                    `P@ףp=
�?             4@p       s                   �k@�}�+r��?             3@q       r                   pj@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?w       x                   �x@�IєX�?             1@������������������������       �        
             0@������������������������       �                     �?z       {                   pb@"pc�
�?             &@������������������������       �                     @|       }                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     @       �                    �?Dc}h��?%             L@�       �                   `a@v�2t5�?            �D@�       �                   �b@�ՙ/�?             5@�       �                   �g@��.k���?             1@�       �                   @_@�����H�?             "@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �s@z�G�z�?             4@�       �                   �b@�����H�?             2@�       �                    �?@4և���?
             ,@�       �                   �a@      �?             @�       �                   @m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@�       �                   h@�p�?�             n@�       �                    �?��t���?�            �m@�       �                    �?�7��?0            �S@�       �                    �?`����֜?+            �Q@������������������������       �        '             O@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                    b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �d@��G�?e            �c@�       �                    �?��[�8��?b             c@�       �       	          ����?����Q8�?.            �Q@�       �                   �a@P����?&            �M@�       �                   �\@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                    �F@�       �                   l@      �?             (@������������������������       �                     @�       �       	          `ff�?      �?             @�       �                    �?      �?             @������������������������       �                     �?�       �                   xp@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @H�U?B�?4            �T@�       �                   @[@���!pc�?&            �K@������������������������       �                     @�       �       	          `ff�?�θ�?%             J@�       �                   `a@Jm_!'1�?#            �H@������������������������       �        	             &@�       �                     H@�I�w�"�?             C@������������������������       �                     0@�       �                     N@8�A�0��?             6@�       �                   �b@     ��?             0@������������������������       �                     @�       �                   �l@�z�G��?             $@������������������������       �                     @�       �       	          ����?      �?             @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     I@|��?���?             ;@�       �                   �l@ףp=
�?             $@�       �                   `f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �p@�t����?	             1@�       �                   �`@$�q-�?             *@�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �                    a@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �h@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          033@ףp=
�?             >@������������������������       �        
             ,@�       �                    �G@     ��?             0@�       �                   (p@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?$�q-�?             *@������������������������       �                     &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�        t@     �y@      M@     p@      G@      N@      7@       @      "@              ,@       @              @      ,@       @      (@               @       @               @       @              7@      J@      @     �@@              $@      @      7@      @              @      7@      @      .@      @      @       @              �?      @      �?                      @              (@               @      1@      3@      0@      "@      .@      @      @      @       @      @              @       @              @              $@              �?      @      �?      �?      �?                      �?              @      �?      $@      �?       @      �?      �?              �?      �?                      �?               @      (@     �h@      "@     @Q@      "@      L@      @      �?      @                      �?      @     �K@       @      I@             �D@       @      "@               @       @      �?              �?       @              @      @              @      @      �?      @                      �?              *@      @      `@       @      `@              Y@       @      <@      �?      �?      �?                      �?      �?      ;@      �?      @      �?                      @              8@      �?             �p@     `c@     Pp@      `@     @P@     �T@      @      4@       @      4@      �?      4@              &@      �?      "@      �?      @               @      �?      �?      �?                      �?              @      �?              �?              O@     �O@     �F@      8@     �E@      .@      ;@      ,@              @      ;@      "@      "@      @      @              @      @              @      @       @               @      @              2@      @      2@       @      2@      �?       @      �?       @                      �?      $@                      �?              �?      0@      �?      0@                      �?       @      "@              @       @      @       @                      @      1@     �C@      1@      8@      *@       @      "@       @       @      �?      @              �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?      @              @      0@       @      0@      �?      *@      �?      @      �?      �?              �?      �?                       @              $@      �?      @              @      �?               @                      .@     �h@     �F@     `h@      E@     �R@      @     @Q@      �?      O@              @      �?              �?      @              @      @      @              �?      @              @      �?             @^@      C@      ^@     �@@     �P@      @      M@      �?      *@      �?              �?      *@             �F@              "@      @      @              @      @      �?      @              �?      �?       @               @      �?               @             �J@      =@      D@      .@              @      D@      (@      D@      "@      &@              =@      "@      0@              *@      "@      @      "@              @      @      @      @              �?      @      �?      �?              �?      �?                       @      @                      @      *@      ,@      �?      "@      �?      @      �?                      @              @      (@      @      (@      �?       @      �?              �?       @              $@                      @      �?      @      �?                      @      �?      @              @      �?              @      ;@              ,@      @      *@       @      �?       @                      �?      �?      (@              &@      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B88         �                    �?0����?�           ��@       A                    �?���\�?�            �x@                          @_@�E��
��?\            �c@                           �?�{��?��?"             K@������������������������       �                      @                           �?D>�Q�?              J@                          �Q@$�q-�?            �C@������������������������       �                      @	                           V@�?�|�?            �B@
              	          ����?���N8�?             5@              	          ���ܿ��S�ۿ?             .@������������������������       �                     @                          �Z@�C��2(�?             &@������������������������       �                     "@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             0@                            P@��
ц��?             *@                           �?���Q��?	             $@                           @L@؇���X�?             @                          `Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @       >                   �b@Np�����?:            �Y@       =                    �?��
ц��?5            �V@       2                   �n@~�hP��?,            �R@        +                   �c@z�G�z�?             D@!       "                    �?�X����?             6@������������������������       �                      @#       *       	          @33�?      �?             4@$       )                   �g@r�q��?             2@%       (                   @_@և���X�?             @&       '                    b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �                      @,       -       	             �?�X�<ݺ?             2@������������������������       �                     (@.       /                     I@r�q��?             @������������������������       �                     @0       1       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?3       <                   �r@      �?             A@4       7                    �?��+7��?             7@5       6                   Pp@�q�q�?             @������������������������       �                      @������������������������       �                     �?8       ;                   @b@z�G�z�?             4@9       :                     N@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@������������������������       �                     &@������������������������       �        	             1@?       @                   �a@���!pc�?             &@������������������������       �                     @������������������������       �                      @B       �                    �N@�����H�?�            `n@C       f                    �?��y�S��?x             h@D       S                    �I@ףp=
�?^            �b@E       R                   �e@ZՏ�m|�?!            �H@F       G                   �Z@��E�B��?             �G@������������������������       �                      @H       K                    �?�:�^���?            �F@I       J       	          ����?      �?             @������������������������       �                      @������������������������       �                      @L       Q       	          `ff�?������?            �D@M       N                    @G@      �?              @������������������������       �                     @O       P                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �@@������������������������       �                      @T       U                    �?�L�L��?=            @Y@������������������������       �                    �A@V       a                   @m@��IF�E�?+            �P@W       `                   `l@     ��?             @@X       Y                    �?�r����?             >@������������������������       �                     �?Z       _                   �`@ܷ��?��?             =@[       \                   �^@�θ�?	             *@������������������������       �                      @]       ^                   �j@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@������������������������       �                      @b       c                    @M@г�wY;�?             A@������������������������       �                     ?@d       e                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?g       t                    @M@�%^�?            �E@h       s                    �?؇���X�?             <@i       p       	             @z�G�z�?             4@j       k                   �[@r�q��?             2@������������������������       �                      @l       o                   �X@      �?
             0@m       n                   @^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@q       r       	             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @u       x                    �?��S���?             .@v       w                   �s@���Q��?             @������������������������       �                      @������������������������       �                     @y       |                    �M@      �?             $@z       {                    _@z�G�z�?             @������������������������       �                     �?������������������������       �                     @}       �                   �a@z�G�z�?             @~                          �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �R@p���?              I@������������������������       �                     H@�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          pff�?V~b���?�            �t@�       �                    I@J�:�Ȣ�?�            �o@�       �                   `_@      �?             0@�       �                    �?ףp=
�?             $@�       �                    `R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    a@r�q��?             @������������������������       �                     @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @��w\ud�?�            �m@�       �                    ]@�Cc}h��?�             l@�       �                   �Z@ �o_��?             9@������������������������       �                     @�       �                   `l@b�2�tk�?             2@������������������������       �                     @�       �                    �?���|���?             &@������������������������       �                     �?�       �                    �?�z�G��?             $@������������������������       �                     @�       �                    �D@      �?             @������������������������       �                      @�       �                   @[@      �?             @������������������������       �                      @�       �                     J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �? l����?}            �h@�       �                   �j@H�_�r�?n            `f@������������������������       �        '            �P@�       �                    �?4�0_���?G            @\@�       �                   �^@ >�֕�?A            @Z@������������������������       �                    �C@�       �                    �?�C��2(�?,            �P@�       �       	            �?�(\����?             D@������������������������       �                    �A@�       �                    _@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   @o@���B���?             :@�       �                     G@���Q��?             $@������������������������       �                     @�       �                     M@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `a@      �?             0@������������������������       �                     $@�       �       	          @33�?r�q��?             @�       �                   �t@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   pb@      �?              @�       �                   �`@      �?             @������������������������       �                      @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �]@�z�G��?             4@������������������������       �                     @�       �                   �`@      �?             0@������������������������       �                      @�       �                   `a@      �?              @������������������������       �                     @�       �                   Pc@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @N@      �?
             ,@�       �                    �?���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ���@^�JB=�?<            @T@�       �                   �d@�9mf��?,            �O@�       �                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                    �?��e�B��?%            �I@�       �                    �?#z�i��?            �D@�       �                    �?$�q-�?             *@������������������������       �                     @�       �                   `o@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �b@���>4��?             <@�       �                    a@����X�?
             ,@�       �                    @X�<ݚ�?             "@�       �                   @m@z�G�z�?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   0e@d}h���?	             ,@�       �                    �?�8��8��?             (@�       �                    p@r�q��?             @������������������������       �                     @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �I@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �?�����H�?             2@������������������������       �                     �?�       �                    �?�IєX�?             1@������������������������       �                     *@�       �                    �?      �?             @������������������������       �                     �?�                           �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�b��     h�h(h+K ��h-��R�(KMKK��h^�B        u@     �x@     �V@     Ps@     �O@     @W@      &@     �E@       @              "@     �E@      @      B@       @              �?      B@      �?      4@      �?      ,@              @      �?      $@              "@      �?      �?              �?      �?                      @              0@      @      @      @      @      @      �?       @      �?              �?       @              @                      @              @      J@      I@     �H@      E@     �H@      9@      @@       @      .@      @               @      .@      @      .@      @      @      @       @      @       @                      @       @              &@                       @      1@      �?      (@              @      �?      @              �?      �?              �?      �?              1@      1@      @      1@       @      �?       @                      �?      @      0@      @       @      @                       @              ,@      &@                      1@      @       @      @                       @      ;@      k@      :@     �d@      .@     �`@       @     �D@      @     �D@       @              @     �D@       @       @       @                       @       @     �C@       @      @              @       @      �?              �?       @                     �@@       @              @     �W@             �A@      @     �M@      @      :@      @      :@      �?              @      :@      @      $@               @      @       @      @                       @              0@       @              �?     �@@              ?@      �?       @               @      �?              &@      @@      @      8@      @      0@      @      .@       @              �?      .@      �?       @               @      �?                      *@      �?      �?      �?                      �?               @      @       @       @      @       @                      @      @      @      @      �?              �?      @              �?      @      �?      �?              �?      �?                      @      �?     �H@              H@      �?      �?      �?                      �?     �n@     @V@     �j@     �C@      @      $@      �?      "@      �?       @               @      �?                      @      @      �?      @              �?      �?      �?                      �?      j@      =@     @i@      6@      2@      @      @              &@      @      @              @      @      �?              @      @              @      @      @       @              �?      @               @      �?      �?              �?      �?              g@      .@     @e@      "@     �P@              Z@      "@     �X@      @     �C@              N@      @     �C@      �?     �A@              @      �?              �?      @              5@      @      @      @      @              �?      @              @      �?              .@      �?      $@              @      �?      @      �?      @                      �?       @              @      @      �?      @               @      �?      �?      �?                      �?      @              ,@      @              @      ,@       @       @              @       @      @               @       @               @       @              @      @      @      @      @                      @      @              ?@      I@      =@      A@      �?      &@      �?                      &@      <@      7@      ;@      ,@      (@      �?      @              @      �?      @               @      �?       @                      �?      .@      *@      @      $@      @      @      �?      @      �?      �?              �?      �?                      @      @      �?              �?      @                      @      &@      @      &@      �?      @      �?      @              �?      �?              �?      �?              @                       @      �?      "@      �?                      "@       @      0@      �?              �?      0@              *@      �?      @              �?      �?       @      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KKᅔh}�B81         l                   �`@�+	G�?�           ��@       Y                    �?l�"�^%�?�            �u@       .       	          ����?0�	B��?�            �n@       )                   `_@D�n�3�?;            �W@                            J@��(@��?-            �Q@                           �?      �?             4@                          �^@X�<ݚ�?             "@������������������������       �                     @	                           @H@�q�q�?             @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@       "                   �k@��H�}�?!             I@                          `c@�s��:��?             C@                           �?��<b���?             7@������������������������       �                     *@                           �?      �?             $@                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?և���X�?             @                          �]@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                           �L@z�G�z�?
             .@������������������������       �                     @       !                    @M@�q�q�?             "@                           @Z@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @#       $                    �?�8��8��?             (@������������������������       �                     "@%       (                   @_@�q�q�?             @&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?*       -                    �?H%u��?             9@+       ,                   �]@�nkK�?             7@������������������������       �                     �?������������������������       �                     6@������������������������       �                      @/       8                    �?h�˹�?g             c@0       1                    i@�����?             3@������������������������       �                      @2       7                    @������?
             1@3       4                   �]@@4և���?             ,@������������������������       �                     &@5       6                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @9       L                    �?ՀJ��?[            �`@:       A                    @M@io8�?N             ]@;       <       	          033@�(�Tw�?3            �S@������������������������       �        +             Q@=       >                    �?ףp=
�?             $@������������������������       �                      @?       @                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?B       K                    �O@�S����?             C@C       H                   P`@����X�?             5@D       G       	          ����?      �?             0@E       F                    @O@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @I       J                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@M       N                     I@�t����?             1@������������������������       �                     @O       X                    @�n_Y�K�?
             *@P       W                    c@�q�q�?	             (@Q       R                   �o@���!pc�?             &@������������������������       �                     @S       T                   �q@���Q��?             @������������������������       �                      @U       V                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?Z       _                    �?�C��2(�?A            �X@[       \                   �b@�q�q�?             "@������������������������       �                     @]       ^                    �?      �?             @������������������������       �                     @������������������������       �                     �?`       a                   �k@��S�ۿ?<            �V@������������������������       �        '             L@b       c                    @G@@�0�!��?             A@������������������������       �                      @d       g                   pm@      �?             @@e       f                    �P@      �?             @������������������������       �                      @������������������������       �                      @h       i                   �S@@4և���?             <@������������������������       �                     �?j       k                    �R@ 7���B�?             ;@������������������������       �                     :@������������������������       �                     �?m       �                    �?�E���?�            @x@n       s                   @E@��ʫf_�?�            �r@o       p                    �N@���N8�?             5@������������������������       �                     3@q       r                    �?      �?              @������������������������       �                     �?������������������������       �                     �?t       �                    �?2L�����?�            @q@u       z                    �?��W3�?*            �Q@v       w                   �b@PN��T'�?             ;@������������������������       �                     6@x       y                   0d@z�G�z�?             @������������������������       �                     @������������������������       �                     �?{       �                    �L@d�
��?             F@|       �       	          ����?�LQ�1	�?             7@}       �                   �d@���!pc�?             &@~       �                    e@�����H�?             "@       �                     F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     (@�       �                   �l@؇���X�?             5@�       �       	          033@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@�       �                   ht@6��m�?�            �i@�       �       	          `ff@�DÓ ��?�            @i@�       �                   �]@(l58��?            �h@�       �                   �a@��R[s�?            �A@������������������������       �                     @�       �                    f@�חF�P�?             ?@�       �                    �?�GN�z�?             6@������������������������       �                     "@�       �                   pd@�n_Y�K�?
             *@�       �                     D@z�G�z�?             $@������������������������       �                     �?�       �                   �n@�����H�?             "@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    @������?h            �d@�       �                    �?`-�I�w�?a             c@�       �                    f@ �Cc}�?             <@�       �                     N@�8��8��?             8@�       �                   �_@���N8�?             5@�       �                   pk@r�q��?             @�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        
             .@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �f@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	            �?�&/�E�?O             _@�       �                    �?@��8��??             X@�       �                    �?��f�{��?8            �U@������������������������       �        2             S@�       �                    �G@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �       	          ����?ףp=
�?             $@�       �                   �b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�>4և��?             <@�       �                    _@��<b���?             7@�       �                   �^@���Q��?             @�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �b@�����H�?	             2@�       �                   �f@�IєX�?             1@������������������������       �                     �?������������������������       �                     0@������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?             (@������������������������       �                     @�       �                    �?      �?              @�       �                     P@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@�DC��,�?2            �V@�       �                   �\@ 	��p�?!             M@�       �                   �m@���Q��?             $@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     H@�       �       	          ����?4���C�?            �@@�       �                    �?�<ݚ�?	             2@������������������������       �                     $@�       �                   �p@      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             .@�       �                   �p@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B       `t@     �y@     �T@     �p@     @R@     �e@     �K@      D@     �@@     �B@      .@      @      @      @              @      @       @      �?       @      �?                       @      @              &@              2@      @@      1@      5@      @      2@              *@      @      @       @      �?              �?       @              @      @      @       @      @                       @               @      (@      @      @              @      @       @      @       @                      @      @              �?      &@              "@      �?       @      �?      �?      �?                      �?              �?      6@      @      6@      �?              �?      6@                       @      2@     �`@      @      *@       @              @      *@      �?      *@              &@      �?       @      �?                       @      @              (@     @^@      @     @[@      �?     @S@              Q@      �?      "@               @      �?      �?      �?                      �?      @      @@      @      .@       @      ,@       @      @              @       @                      @      @      �?              �?      @                      1@      @      (@              @      @       @      @       @      @       @              @      @       @       @              �?       @      �?                       @      �?              �?              "@     �V@      @      @              @      @      �?      @                      �?      @      U@              L@      @      <@       @              @      <@       @       @               @       @               @      :@      �?              �?      :@              :@      �?             �n@      b@     �k@      S@      �?      4@              3@      �?      �?              �?      �?             �k@      L@      G@      9@      7@      @      6@              �?      @              @      �?              7@      5@      4@      @       @      @       @      �?       @      �?              �?       @              @                       @      (@              @      2@      @       @      @                       @              0@     �e@      ?@     �e@      <@     �e@      9@      :@      "@              @      :@      @      1@      @      "@               @      @       @       @              �?       @      �?      @      �?      @                      �?      @                      @      "@             �b@      0@     �a@      $@      9@      @      6@       @      4@      �?      @      �?       @      �?       @                      �?      @              .@               @      �?       @                      �?      @      �?              �?      @             @]@      @     �W@       @     @U@      �?      S@              "@      �?              �?      "@              "@      �?      @      �?              �?      @              @              7@      @      2@      @       @      @       @      �?              �?       @                       @      0@       @      0@      �?              �?      0@                      �?      @              @      @      @               @      @      �?      @              @      �?              �?                      @              @      7@      Q@      @      K@      @      @      @      �?              �?      @                      @              H@      3@      ,@      ,@      @      $@              @      @      @                      @      @      $@       @      $@              $@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK�h}�B(5         �                    �?6������?�           ��@                           �?(��3Ea�?�             w@                          �R@N1���?'            �N@������������������������       �                     "@                           �J@��
ц��?!             J@                          `c@z�G�z�?             9@              	          ����?r�q��?             8@������������������������       �        
             3@	       
                   �`@z�G�z�?             @������������������������       �                     @                          Pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           �P@l��
I��?             ;@              	          ����?�㙢�c�?             7@              	          @33�?X�<ݚ�?             "@������������������������       �                     @                            P@�q�q�?             @                           �?z�G�z�?             @                           �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        	             ,@������������������������       �                     @       [                    �?N��s�?�            0s@       N       	          ����?�{���2�?M            �[@       A                   ``@P��E��?/             R@       <                    �?�q����?#            �J@        ;                    @O@��]�T��?            �D@!       :                   �f@��Q��?             D@"       9                    �?�����?             C@#       8                   po@��R[s�?            �A@$       7                   �k@�q�q�?             ;@%       6       	             �? �o_��?             9@&       -                   `Z@�q�q�?             8@'       ,                   @E@և���X�?             @(       )                   �_@���Q��?             @������������������������       �                      @*       +                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @.       /                   �h@@�0�!��?             1@������������������������       �                     "@0       3                    �?      �?              @1       2                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?4       5                   �b@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?=       >                   �l@�8��8��?             (@������������������������       �                     "@?       @       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?B       K                    �?�����?             3@C       J       	             �?X�Cc�?             ,@D       E                     E@�q�q�?             (@������������������������       �                      @F       I                    m@�z�G��?             $@G       H                   �^@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @L       M                    @P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?O       Z                   �t@�ݜ�?            �C@P       Y                    �?�L���?            �B@Q       R                   �U@؇���X�?             5@������������������������       �                      @S       X                    @K@�}�+r��?             3@T       U                    �J@�����H�?             "@������������������������       �                     @V       W                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     0@������������������������       �                      @\       �                   �d@Hm_!'1�?�            �h@]       �                    �R@�v�|�<�?            �g@^       _                   �U@8v�YeK�?~            �g@������������������������       �                      @`       �                   0c@��ɹ?}            �g@a       �                   0c@x��-�?j            �c@b       �                   Hq@Х-��ٹ?d            �b@c       d                    �F@T(y2��?O            �]@������������������������       �                     6@e       p       	          hff�?DE�SA_�?B            @X@f       o                   �b@      �?             0@g       h                   �_@؇���X�?             ,@������������������������       �                      @i       n                   �^@�q�q�?             @j       k                    �O@z�G�z�?             @������������������������       �                     @l       m                   0o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q       z                   @l@H�!b	�?6            @T@r       s                    �M@ pƵHP�?#             J@������������������������       �                    �@@t       u       	          ����?�}�+r��?             3@������������������������       �                     &@v       y       	             @      �?              @w       x                   @`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @{       �                    �?ܷ��?��?             =@|                           @G@ �Cc}�?             <@}       ~       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `\@$�q-�?             :@�       �                   `[@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �        
             0@������������������������       �                     �?������������������������       �                     ?@�       �                   �p@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     =@������������������������       �                     �?�       �                   Pe@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?H��Ly��?�            �v@�       �       	          ���@��11��?�            �r@�       �                   Hp@T;���?�            �q@�       �                   �c@�P�U`��?�            `h@�       �       	          ����?�G��l��?             5@�       �                    @���!pc�?             &@�       �                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �_@z�G�z�?             $@�       �                   `^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�8���?y            �e@������������������������       �        <            @T@�       �                    Z@��a�n`�?=            @W@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @L@����\�?:            �V@�       �                   Pd@      �?,             P@������������������������       �                     A@�       �                   �n@��S�ۿ?             >@�       �                   m@h�����?             <@������������������������       �                     6@�       �                   @m@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?���B���?             :@�       �                    d@      �?             8@�       �                   �l@�IєX�?	             1@������������������������       �                     &@�       �                   �l@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	          033�?����X�?             @�       �                   �i@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?Z��:���?1            �V@�       �       	          ����?HP�s��?             9@������������������������       �                     3@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?8�A�0��?             �P@�       �                   �d@�-ῃ�?            �N@�       �                    d@�����?            �L@�       �       	          ����?�xGZ���?            �A@�       �                    @��X��?             <@�       �                   Pa@�㙢�c�?             7@������������������������       �                     $@�       �       	          ����?�	j*D�?             *@�       �                   �c@���Q��?             $@�       �                    �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   `]@�C��2(�?             6@������������������������       �                      @������������������������       �                     4@������������������������       �                     @������������������������       �                     @�       �                   �i@$�q-�?	             *@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �b@P�~D&�?+            �P@�       �                   �r@PN��T'�?#             K@�       �                    �J@�8��8��?             H@�       �                    �?�θ�?             *@������������������������       �                      @�       �                    `@�C��2(�?             &@������������������������       �                      @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?��?^�k�?            �A@�       �                    _@@4և���?             ,@������������������������       �                     &@�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     5@�       �                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �C@�θ�?             *@������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h^�B0       �t@     �x@     �S@      r@      <@     �@@              "@      <@      8@      4@      @      4@      @      3@              �?      @              @      �?      �?      �?                      �?              �?       @      3@      @      3@      @      @              @      @       @      @      �?      �?      �?              �?      �?              @                      �?              ,@      @              I@     p@      A@     @S@      =@     �E@      0@     �B@      .@      :@      ,@      :@      (@      :@      "@      :@      "@      2@      @      2@      @      1@      @      @       @      @               @       @      �?       @                      �?       @              @      ,@              "@      @      @      �?      �?      �?                      �?       @      @              @       @                      �?       @                       @      @               @              �?              �?      &@              "@      �?       @               @      �?              *@      @      "@      @      @      @               @      @      @      @      @              @      @              @               @              @      �?      @                      �?      @      A@      @      A@      @      2@       @              �?      2@      �?       @              @      �?       @               @      �?                      $@              0@       @              0@     �f@      *@     @f@      (@     @f@       @              $@     @f@      $@     �b@       @     �a@       @     �[@              6@       @     @V@      @      (@       @      (@               @       @      @      �?      @              @      �?      �?              �?      �?              �?               @              @     @S@      �?     �I@             �@@      �?      2@              &@      �?      @      �?      @      �?                      @              @      @      :@      @      9@      �?      �?      �?                      �?       @      8@       @       @               @       @                      0@              �?              ?@       @      @              @       @                      =@      �?              @       @      @                       @     p@     @[@     �m@      N@     �m@      H@      f@      3@      &@      $@      @       @      @       @               @      @                      @       @       @       @       @       @                       @      @             �d@      "@     @T@              U@      "@      �?       @      �?                       @     �T@      @      O@       @      A@              <@       @      ;@      �?      6@              @      �?              �?      @              �?      �?              �?      �?              5@      @      5@      @      0@      �?      &@              @      �?              �?      @              @       @       @       @               @       @              @                       @      O@      =@      7@       @      3@              @       @               @      @             �C@      ;@     �C@      6@     �C@      2@      3@      0@      3@      "@      3@      @      $@              "@      @      @      @      �?      @      �?                      @      @              @                      @              @      4@       @               @      4@                      @              @      �?      (@               @      �?      @      �?                      @      2@     �H@       @      G@      @      F@      @      $@       @              �?      $@               @      �?       @      �?                       @      �?      A@      �?      *@              &@      �?       @      �?                       @              5@      @       @      @                       @      $@      @              @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK���h}�B�7         �                    �?�Z���?�           ��@                          �`@~�Q7:�?           �z@                           �?O�o9%�?0            �Q@                           �?
j*D>�?             :@������������������������       �                     @              	          �����
;&����?             7@������������������������       �                     @                          �`@�q�q�?             2@	       
                   �Z@�t����?             1@������������������������       �                     @                           �?�n_Y�K�?	             *@                          �[@      �?              @������������������������       �                     �?                          �`@؇���X�?             @������������������������       �                     @                          @E@      �?              @������������������������       �                     �?������������������������       �                     �?                            @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?                          �c@`Ӹ����?            �F@������������������������       �                     A@              	          `ff@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @       }       	          033�?^;|��?�            Pv@       X                    @L@vAƠB��?�            `t@       ;                    �?�J�4�?�             l@       (                   �`@���>4��?#             L@        !                   0g@�t����?             1@������������������������       �                     �?"       #                    �?      �?
             0@������������������������       �                     @$       %                   @_@$�q-�?             *@������������������������       �                     @&       '                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?)       .                   �b@�99lMt�?            �C@*       +                   �`@��S�ۿ?	             .@������������������������       �                     (@,       -                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @/       :                   @t@r�q��?             8@0       3                   @c@�ՙ/�?             5@1       2                   `e@؇���X�?             @������������������������       �                     �?������������������������       �                     @4       7                   �d@      �?             ,@5       6                   `i@؇���X�?             @������������������������       �                     �?������������������������       �                     @8       9       	             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @<       W                    �? 
��р�?o             e@=       @                   �c@x��-�?j            �c@>       ?                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?A       V                   h@0G���ջ?h            �c@B       G                    ]@��F��?g            `c@C       D                   @m@     ��?             0@������������������������       �                     "@E       F                    �I@և���X�?             @������������������������       �                     @������������������������       �                     @H       I                   Pc@~t�8��?Z            `a@������������������������       �        *            �P@J       O       	          ����?���;QU�?0            @R@K       N                   pc@ �Jj�G�?%            �K@L       M                     @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        !             I@P       U                   Pm@�<ݚ�?             2@Q       R                   �c@և���X�?             @������������������������       �                      @S       T       	          pff�?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     &@������������������������       �                     �?������������������������       �                     $@Y       x                    �?���!x��?:            @Y@Z       a                    �?�c�Α�?0            �U@[       \       	          `ff�?      �?             @@������������������������       �                     5@]       `                    �?"pc�
�?             &@^       _       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @b       c                   �h@���Q��?            �K@������������������������       �                     $@d       e                   j@�ݏ^���?            �F@������������������������       �                     @f       i                   �\@\�Uo��?             C@g       h                   @Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @j       w                   �q@�q�q�?            �@@k       l                   �n@>���Rp�?             =@������������������������       �                     $@m       n                   �p@p�ݯ��?             3@������������������������       �                     @o       p                    q@z�G�z�?             .@������������������������       �                     @q       v                   �b@�q�q�?             "@r       s                   �]@؇���X�?             @������������������������       �                     @t       u                    �N@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @y       |                   `c@����X�?
             ,@z       {                    �M@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @~                           ^@r֛w���?             ?@������������������������       �                      @�       �                    �?V�a�� �?             =@�       �                   �o@H%u��?             9@�       �                   Pm@      �?             (@�       �       	          033�?�����H�?	             "@������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?$��n�?�             s@�       �                    �?؇���X�?�            �m@�       �                    `@�E5;5 �?t            �e@�       �                    \@d/
k�?H             [@�       �                   Hs@Riv����?$             M@�       �                   �k@ףp=
�?!             I@�       �                    @L@(;L]n�?             >@������������������������       �        	             1@�       �                   �X@$�q-�?
             *@�       �                    @M@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �p@z�G�z�?             4@�       �                   �`@X�<ݚ�?             "@�       �                   �^@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    Z@      �?              @������������������������       �                     @������������������������       �                     @�       �                    @L@`2U0*��?$             I@������������������������       �                     <@�       �                    _@�C��2(�?             6@�       �       	          ����?���N8�?             5@�       �                    �N@ףp=
�?             $@�       �                     N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     �?�       �       	          ����?�%o��?,            �P@�       �       	          033�?�ՙ/�?             E@�       �                    �F@����X�?            �A@������������������������       �                     @�       �                    f@�q�q�?             >@�       �                   �[@�θ�?             :@�       �                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   pm@؇���X�?             5@�       �                    �?      �?             @������������������������       �                      @�       �                     M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             .@������������������������       �                     @�       �                   �`@؇���X�?             @������������������������       �                     @�       �                    Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?z�G�z�?             9@������������������������       �                     �?�       �                   �a@�q�q�?             8@������������������������       �        	             *@�       �                     K@�eP*L��?             &@�       �                    \@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       	             @z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �p@�i�y�?(            �O@������������������������       �                     H@�       �                   `_@�r����?
             .@�       �                   0r@�q�q�?             @������������������������       �                     �?�       �                    �Q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                    I@<��¤�?,             Q@�       �       	          ����?�t����?             1@������������������������       �                     "@�       �                    �?      �?              @�       �                    �M@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    �?Np�����?!            �I@�       �                   �b@      �?             D@�       �                    �?<ݚ)�?             B@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                   @`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     N@���Q��?             9@�       �       	             �?�z�G��?             4@�       �                    ]@      �?             0@������������������������       �                     @�       �                   �b@���Q��?             $@�       �                   �r@      �?              @�       �                    �K@؇���X�?             @������������������������       �                     @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    a@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�        u@     �x@     Pq@     �b@      *@      M@      &@      .@              @      &@      (@      @              @      (@      @      (@              @      @       @       @      @      �?              �?      @              @      �?      �?              �?      �?              @       @      @                       @      �?               @     �E@              A@       @      "@              "@       @             �p@     @W@      p@     �Q@     �g@      B@      >@      :@      @      (@      �?              @      (@      @              �?      (@              @      �?      @              @      �?              9@      ,@      ,@      �?      (@               @      �?              �?       @              &@      *@       @      *@      �?      @      �?                      @      @      @      @      �?              �?      @              �?      @              @      �?              @             �c@      $@     �b@      $@       @      �?       @                      �?     `b@      "@     `b@       @      *@      @      "@              @      @              @      @             �`@      @     �P@              Q@      @      K@      �?      @      �?      @                      �?      I@              ,@      @      @      @               @      @       @               @      @              &@                      �?      $@             �P@      A@     �O@      8@      >@       @      5@              "@       @      @       @               @      @              @             �@@      6@      $@              7@      6@              @      7@      .@      �?      @      �?                      @      6@      &@      6@      @      $@              (@      @              @      (@      @      @              @      @      @      �?      @              @      �?      @                      �?               @              @      @      $@      @      @      @                      @              @       @      7@       @              @      7@      @      6@      @      "@      �?       @      �?                       @       @      �?              �?       @                      *@      @      �?              �?      @             �N@     �n@      A@     �i@      @@     �a@      &@     @X@      "@     �H@      @     �F@      �?      =@              1@      �?      (@      �?      @      �?                      @              @      @      0@      @      @      @      �?              �?      @              �?      @      �?      �?      �?                      �?              @              &@      @      @              @      @               @      H@              <@       @      4@      �?      4@      �?      "@      �?      @              @      �?                      @              &@      �?              5@      G@      0@      :@      $@      9@              @      $@      4@      @      4@      @       @      @                       @      @      2@      @      @               @      @      �?      @                      �?              .@      @              @      �?      @               @      �?       @                      �?      @      4@              �?      @      3@              *@      @      @      @       @      @                       @      �?      @      �?                      @       @     �N@              H@       @      *@       @      @      �?              �?      @              @      �?                      "@      ;@     �D@       @      .@              "@       @      @       @      @              @       @                      �?      9@      :@      9@      .@      9@      &@      $@      �?      @              @      �?              �?      @              .@      $@      ,@      @      $@      @      @              @      @       @      @      �?      @              @      �?      �?              �?      �?              �?               @              @              �?      @      �?                      @              @              &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuMhvh(h+K ��h-��R�(KM��h}�B�8         t                   �`@�#i����?�           ��@       =                    �?����m�?�            �r@       "                    �?���Q��?M            �[@       !                   �e@���}D�?,            �P@                          �\@     ��?+             P@                           �?      �?	             0@������������������������       �                     @       	                    [@r�q��?             (@������������������������       �                      @
              	          `ff�?      �?             @                           �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                            �?8��8���?"             H@                          �k@ �o_��?             9@                           �?p�ݯ��?             3@              	             �?d}h���?             ,@                          �V@      �?             @������������������������       �                     �?                          �O@���Q��?             @������������������������       �                     �?                          �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           `@z�G�z�?             @������������������������       �                      @                           @J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     7@������������������������       �                     @#       2                   �a@8�$�>�?!            �E@$       )                   �\@�q�q�?             8@%       (                    @      �?             @&       '                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @*       /       	             �?ףp=
�?             4@+       .                   @V@�X�<ݺ?             2@,       -                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@0       1                   @[@      �?              @������������������������       �                     �?������������������������       �                     �?3       :                    �?�\��N��?             3@4       5                    �?�z�G��?             $@������������������������       �                      @6       9                     Q@      �?              @7       8                    @L@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @;       <                    �L@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @>       S                   Pl@x�����?~            �g@?       F                    �?�h����?K             \@@       E                   �[@ Df@��?7            �T@A       B                    Y@      �?             0@������������������������       �                     (@C       D                   pi@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        /            �P@G       R                    �?\-��p�?             =@H       O                   �b@      �?             0@I       N       	          033�?�8��8��?             (@J       M                    a@r�q��?             @K       L                   �X@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @P       Q                    �N@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             *@T       W                   �l@��t���?3            �S@U       V                   @`@      �?             @������������������������       �                     �?������������������������       �                     @X       i                    �?���?0            �R@Y       d                   ``@     p�?(             P@Z       [                   �_@�㙢�c�?             7@������������������������       �                     .@\       ]                   Pp@      �?              @������������������������       �                      @^       c                    �?�q�q�?             @_       b                    �?z�G�z�?             @`       a                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?e       f                    �?��Y��]�?            �D@������������������������       �                     @@g       h                    �I@�����H�?             "@������������������������       �                     �?������������������������       �                      @j       s       	          @33�?�eP*L��?             &@k       p                    �?���Q��?             $@l       m                    �?���Q��?             @������������������������       �                     �?n       o                    d@      �?             @������������������������       �                      @������������������������       �                      @q       r                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?u       �                    �?F�Q�j�?           {@v       �       	          ��� @V~b���?�            �t@w       |                   �O@�<ݚ�?�            �s@x       {                    �?`2U0*��?             9@y       z                   @_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@}       �                    �?<�&9�?�             r@~                           �?0�>���?4            �V@������������������������       �                     C@�       �                   �g@0��_��?            �J@�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     @�       �                   �`@����?�?            �F@������������������������       �                     =@�       �                    �H@      �?
             0@������������������������       �                     �?������������������������       �        	             .@�       �                    �?�k�>��?y            �h@�       �                    �?4���C�?'            �P@�       �                   pf@�θ�?	             *@������������������������       �                     $@������������������������       �                     @�       �                    �?r�z-��?            �J@�       �       	          ����?      �?             H@�       �                     M@�g�y��?             ?@�       �                   �_@և���X�?             <@�       �                   �^@X�Cc�?	             ,@�       �                   @b@�q�q�?             (@������������������������       �                     @�       �                    �B@�<ݚ�?             "@������������������������       �                     �?�       �                   pi@      �?              @������������������������       �                     @�       �                    �D@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �a@d}h���?	             ,@������������������������       �                     $@�       �                    d@      �?             @������������������������       �                      @�       �                   �s@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    `P@@�0�!��?             1@�       �                   pj@��S�ۿ?             .@������������������������       �                     "@�       �                   �b@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @pJQg���?R            �`@�       �                   �[@0{�v��?K            @_@�       �                   �d@z�G�z�?             4@�       �                   @c@@4և���?             ,@�       �                   @[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                    �?      �?             @�       �       	             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    @L@���N8�?C            @Z@������������������������       �        5            �T@�       �                    @M@��<b���?             7@�       �       	            �?���|���?             &@�       �                   �h@      �?              @������������������������       �                     @�       �                   �k@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �O@�8��8��?             (@������������������������       �                     $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                     @�       �                   `c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?P���Q�?             4@������������������������       �        
             *@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�J��%�?<            �X@�       �                   �b@\X��t�?             7@�       �                    �?$�q-�?
             *@�       �                    @O@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �P@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                    @I@�M;q��?-            �R@�       �       	             �?      �?             0@�       �                   c@r�q��?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �       	              @�z�G��?             $@�       �                   @`@և���X�?             @�       �                    �?���Q��?             @�       �                    �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �a@��mo*�?"            �M@�       �                    �?��.k���?             1@�       �                    �N@"pc�
�?             &@�       �                    �?�q�q�?             @�       �                   �`@���Q��?             @������������������������       �                     �?�       �                    �J@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@؇���X�?             E@������������������������       �                     7@�                          �?�����?	             3@�             	          ����?@4և���?             ,@�                          @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     @�t�b�5     h�h(h+K ��h-��R�(KMKK��h^�B0       `u@     �x@      P@     �m@      F@     �P@      0@     �I@      *@     �I@      @      $@      @               @      $@               @       @       @       @      �?       @                      �?              �?      @     �D@      @      2@      @      (@      @      &@      @      @              �?      @       @      �?               @       @               @       @                       @      @      �?       @               @      �?              �?       @                      @              7@      @              <@      .@      3@      @      �?      @      �?      �?              �?      �?                       @      2@       @      1@      �?       @      �?              �?       @              .@              �?      �?              �?      �?              "@      $@      @      @       @              @      @       @      @       @                      @      @               @      @       @                      @      4@     `e@      @     �Z@       @     @T@       @      ,@              (@       @       @       @                       @             �P@      @      9@      @      (@      �?      &@      �?      @      �?      @      �?                      @              �?              @      @      �?      @                      �?              *@      ,@     @P@      @      �?              �?      @              &@      P@      @     �M@      @      3@              .@      @      @               @      @       @      @      �?       @      �?       @                      �?       @                      �?      �?      D@              @@      �?       @      �?                       @      @      @      @      @       @      @              �?       @       @       @                       @      @      �?              �?      @                      �?     `q@     `c@     �n@     @V@     �n@     �Q@      �?      8@      �?      @              @      �?                      4@     �n@      G@     �U@      @      C@              H@      @      @      @      @                      @      F@      �?      =@              .@      �?              �?      .@             �c@     �D@      C@      <@      @      $@              $@      @             �A@      2@      >@      2@      0@      .@      0@      (@      @      "@      @      @      @               @      @      �?              �?      @              @      �?      @              @      �?                       @      &@      @      $@              �?      @               @      �?      �?              �?      �?                      @      ,@      @      ,@      �?      "@              @      �?              �?      @                       @      @              ^@      *@      ]@      "@      0@      @      *@      �?      @      �?              �?      @              "@              @      @       @      @       @                      @      �?              Y@      @     �T@              2@      @      @      @      @      �?      @              @      �?              �?      @                      @      &@      �?      $@              �?      �?      �?                      �?      @      @              @      @      �?      @                      �?      �?      3@              *@      �?      @              @      �?              @@     �P@      $@      *@      �?      (@      �?      @              @      �?                      @      "@      �?      "@                      �?      6@     �J@       @       @      @      �?      @      �?      @                      �?       @              @      @      @      @      @       @       @       @              �?       @      �?              �?       @              �?                       @              @      ,@     �F@       @      "@       @      "@       @      @       @      @      �?              �?      @      �?                      @              �?              @      @              @      B@              7@      @      *@      �?      *@      �?      �?      �?                      �?              (@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK݅�h}�BX0         0                    �?"��G,�?�           ��@                          �R@� ��fd�?a            @b@                           @O@؇���X�?             @������������������������       �                     @������������������������       �                     �?       /       	          ���@lQ���?Z            `a@                           �?@�0�!��?Y             a@              	          `ff�?�q-�?E             Z@	                           �?h�a��?@            @X@
                           �?���y4F�?             3@                           b@8�Z$���?	             *@������������������������       �                     &@������������������������       �                      @                           �?�q�q�?             @������������������������       �                     @������������������������       �                      @              	          pff�?�(�Tw�?4            �S@������������������������       �        ,             P@                          �p@@4և���?             ,@              	          ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                           �?����X�?             @                            F@�q�q�?             @������������������������       �                     �?                            K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                    �?     ��?             @@        !                   0u@r�q��?             @������������������������       �                     @������������������������       �                     �?#       ,                    �?�n_Y�K�?             :@$       '                   pl@�LQ�1	�?             7@%       &                    `@����X�?             @������������������������       �                      @������������������������       �                     @(       +                   `^@     ��?	             0@)       *                   �Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@-       .                   �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @1       �                    �?V��f_�?]           `�@2       w       	          ����?      �?�            �s@3       P                    �?���P?-�?|            @i@4       5                    T@�q�q�?+            �R@������������������������       �        	             0@6       K                    @N@�Ƀ aA�?"            �M@7       B                   �_@z�J��?            �G@8       A                   �f@�	j*D�?             :@9       :                   �Y@"pc�
�?             6@������������������������       �                     @;       @                   `n@�}�+r��?
             3@<       =                    �?      �?              @������������������������       �                     @>       ?                   �c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @C       J                    �G@���N8�?             5@D       E                   l@      �?             $@������������������������       �                     @F       I                   0a@r�q��?             @G       H                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        	             &@L       O                   @_@�8��8��?             (@M       N                    �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@Q       V                   @[@�i��b��?Q            �_@R       S                    �G@����X�?             @������������������������       �                     @T       U                   �Z@      �?             @������������������������       �                      @������������������������       �                      @W       \                   �c@�r����?N             ^@X       [                    @      �?             @Y       Z                   `Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @]       ^                    X@X�X\,��?H            �\@������������������������       �                     �?_       `                    @H@hdpZ�L�?G            @\@������������������������       �        "             K@a       p                   Hp@$gv&��?%            �M@b       c                    �?�:�^���?            �F@������������������������       �                     6@d       m       	          pff�?�㙢�c�?             7@e       l       	          ����?�KM�]�?             3@f       k                     P@"pc�
�?             &@g       h                    @L@ףp=
�?             $@������������������������       �                     @i       j                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @n       o                   a@      �?             @������������������������       �                      @������������������������       �                      @q       v                    �?և���X�?	             ,@r       s                   xp@�q�q�?             "@������������������������       �                      @t       u                   �d@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @x       �                   �r@�I�w�"�??            �\@y       �                    �?"��3؞�?<            @[@z       �       	          033�?��M���?$             Q@{       �                    �?�'�=z��?            �@@|       }                    �?      �?             (@������������������������       �                     �?~       �       	          033�?���!pc�?             &@       �                   �`@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @�q�q�?             5@�       �                    �?p�ݯ��?             3@�       �                   �\@��S���?	             .@������������������������       �                     @�       �                   @_@�����H�?             "@�       �                   pq@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   pe@ >�֕�?            �A@�       �                   �d@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     :@�       �                   `c@��p\�?            �D@������������������������       �                    �@@�       �       	             @      �?              @�       �                    o@r�q��?             @�       �                    @H@�q�q�?             @������������������������       �                     �?�       �                    @L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �b@`RC4%�?�             q@�       �       	          ����?|�(��?�            �o@�       �                    �D@      �?             J@������������������������       �                     @�       �       	          ����?�����?            �H@�       �                   @a@�����H�?             B@������������������������       �        	             0@�       �                    _@z�G�z�?
             4@�       �                   �T@@4և���?             ,@�       �                    �?؇���X�?             @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                   �i@��
ц��?             *@������������������������       �                     @������������������������       �                     @�       �                    @@,Ԛ��?{             i@�       �                    �?�7f8���?z            �h@�       �                   P`@��X�-�?V            `a@�       �                   `_@�S����?#            �L@�       �                    �?��S�ۿ?             >@�       �                   �^@@4և���?             <@������������������������       �        
             2@�       �                   �_@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �       	          ����?������?             ;@�       �                    `@      �?             $@������������������������       �                     @������������������������       �                     @�       �                    �H@�t����?
             1@�       �                    �D@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @\@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �        3            �T@�       �                   `b@ _�@�Y�?$             M@������������������������       �                     F@�       �       	          ����?@4և���?	             ,@�       �                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @�       �       	          033�?�G�z��?             4@�       �                    @M@�C��2(�?             &@������������������������       �                      @�       �                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �o@�����H�?             "@������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       @s@     �z@     @\@     �@@      �?      @              @      �?              \@      ;@      \@      8@     @X@      @      W@      @      .@      @      &@       @      &@                       @      @       @      @                       @     @S@      �?      P@              *@      �?      @      �?              �?      @              "@              @       @      �?       @              �?      �?      �?      �?                      �?      @              .@      1@      @      �?      @                      �?      $@      0@       @      .@      @       @               @      @              @      *@      @      �?              �?      @                      (@       @      �?       @                      �?              @     `h@     �x@     �c@     �c@     ``@     �Q@      9@      I@              0@      9@      A@      8@      7@       @      2@      @      2@      @              �?      2@      �?      @              @      �?      @              @      �?                      &@      @              0@      @      @      @              @      @      �?       @      �?       @                      �?      @              &@              �?      &@      �?       @      �?                       @              "@     �Z@      5@       @      @              @       @       @       @                       @      Z@      0@      @      @      @      �?              �?      @                       @     @Y@      *@              �?     @Y@      (@      K@             �G@      (@     �D@      @      6@              3@      @      1@       @      "@       @      "@      �?      @              @      �?      @                      �?              �?       @               @       @       @                       @      @       @      @      @               @      @      �?      @                      �?              @      ;@     �U@      6@     �U@      3@     �H@      1@      0@      @      "@              �?      @       @      �?       @               @      �?               @              ,@      @      (@      @       @      @              @       @      �?       @      �?       @                      �?      @              @               @               @     �@@       @      @              @       @                      :@      @      C@             �@@      @      @      �?      @      �?       @              �?      �?      �?      �?                      �?              @       @              @             �B@     `m@      :@     @l@      *@     �C@      @              $@     �C@      @      @@              0@      @      0@      �?      *@      �?      @      �?      @              @      �?                       @              @      @      @              @      @              @      @              @      @              *@     `g@      $@     `g@      "@     @`@      "@      H@       @      <@       @      :@              2@       @       @       @                       @               @      @      4@      @      @      @                      @       @      .@      �?       @               @      �?              �?      *@      �?                      *@             �T@      �?     �L@              F@      �?      *@      �?       @               @      �?                      &@      @              &@      "@      $@      �?       @               @      �?       @                      �?      �?       @              @      �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK���h}�BX7         �       	          ����?�#i����?�           ��@              	          433ӿ`�&�	��?�            �w@������������������������       �                     @       #                   `_@&�
�M�?�            �w@                          b@t�C�#��?7            �S@                          �b@      �?             @@������������������������       �                     8@       	                    �?      �?              @������������������������       �                     @
                          �c@      �?             @������������������������       �                     �?������������������������       �                     @                           �?��C���?            �G@                          �Z@8�A�0��?             6@                          @W@�����H�?             "@������������������������       �                     @              	          ����?z�G�z�?             @                          �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @              	          hff�?$�q-�?	             *@������������������������       �                     &@                            L@      �?              @������������������������       �                     �?������������������������       �                     �?       "                    �?�+e�X�?             9@                           �L@�����?             5@������������������������       �        
             .@                           �?�q�q�?             @������������������������       �                     @        !                    b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @$       s                    �?�w1�|�?�            �r@%       D                   p@�������?�            `p@&       '                    �?���C"��?j            �d@������������������������       �                    �C@(       1                    �?ĭ����?L            @_@)       *                    �D@������?             ;@������������������������       �                     @+       ,                   �b@�LQ�1	�?             7@������������������������       �                     0@-       .                     I@և���X�?             @������������������������       �                     @/       0                   Pk@      �?             @������������������������       �                     @������������������������       �                     �?2       7                    @A@��<D�m�?8            �X@3       4                    �@@�q�q�?             @������������������������       �                     @5       6                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?8       A                    �P@�nkK�?3             W@9       :                   �l@ qP��B�?0            �U@������������������������       �        %             Q@;       <                   �[@�����H�?             2@������������������������       �                     �?=       >                   �`@�IєX�?
             1@������������������������       �                     .@?       @                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?B       C                     Q@�q�q�?             @������������������������       �                      @������������������������       �                     @E       r                    @H��%�R�?7            �X@F       G                   �`@�uw\l��?5            @W@������������������������       �                     @H       g                   pt@>��C��?1            �U@I       R                   �p@z�G�z�?*            �R@J       Q                   �p@b�2�tk�?             2@K       P                   c@     ��?
             0@L       M                    �?����X�?             @������������������������       �                     �?N       O                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @S       \                   �d@Ԫ2��?            �L@T       U                   `b@������?            �D@������������������������       �                     .@V       W                    �C@$�q-�?             :@������������������������       �                     �?X       Y                   �r@`2U0*��?             9@������������������������       �        
             5@Z       [                   s@      �?             @������������������������       �                     �?������������������������       �                     @]       f                   �_@      �?             0@^       e       	             �?�q�q�?             "@_       d                   �^@      �?             @`       a                     C@      �?             @������������������������       �                      @b       c                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @h       i                    �?�eP*L��?             &@������������������������       �                     @j       q                    �?      �?              @k       p                    �N@      �?             @l       o                    �?      �?             @m       n                   8|@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @t       u                    �F@���Q��?            �A@������������������������       �                     @v       �                    �?     ��?             @@w       �       	          ����?�z�G��?             >@x       {                   ``@$��m��?             :@y       z                    �I@r�q��?             @������������������������       �                     �?������������������������       �                     @|       �                    �?z�G�z�?             4@}       ~                   @d@      �?	             0@������������������������       �                     ,@       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?
�GN��?�             v@�       �       	          ���@4���C�?)            �P@�       �       	          ����?l��[B��?$             M@������������������������       �                     @�       �                   �c@�eP*L��?#            �K@�       �                    �?`�(c�?            �H@�       �                    @�q�q�?             2@�       �                    �?      �?	             (@�       �                    �L@      �?              @������������������������       �                     @�       �                    �N@�q�q�?             @������������������������       �                     �?�       �                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?��a�n`�?             ?@�       �       	          ����?8�Z$���?             :@�       �                    �N@�<ݚ�?             2@�       �                   �^@����X�?	             ,@������������������������       �                     @�       �                   @_@�C��2(�?             &@������������������������       �                     @�       �       	          ����?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �K@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   �c@��8���?�            �q@�       �                    _@����a�?�            �n@�       �                    @b�h�d.�?.            �Q@�       �                   pa@��2(&�?+            �P@�       �                    �? �#�Ѵ�?            �E@�       �                    �I@ 	��p�?             =@������������������������       �                     (@�       �                    �J@�t����?             1@������������������������       �                     �?�       �                   `k@      �?             0@�       �                    �?      �?             @�       �                   Ph@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �        	             ,@�       �                    �?8����?             7@�       �                    �H@��S�ۿ?             .@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    @K@      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �e@��-��ĳ?s            �e@�       �       	          ����?���U�?p            `e@�       �                   P`@`Jj��?F            @W@�       �                   �x@x�G�z�?=             T@�       �       	          ����? ���J��?;            �S@�       �                    �? 	��p�?             =@�       �                   �`@ ��WV�?             :@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                   �X@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             0@�       �                   p`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        '            �H@�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   p`@�θ�?	             *@�       �                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �        *            �S@�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    b@      �?             E@�       �                    �?�s��:��?             C@�       �       	             @\X��t�?             7@�       �                     L@������?             1@�       �                    �F@@4և���?
             ,@������������������������       �                     &@�       �                     I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �N@������?             .@�       �                    �?8�Z$���?             *@������������������������       �                     @�       �                    o@����X�?             @�       �                    e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       `u@     �x@      q@      [@              @      q@     �Y@      =@      I@      �?      ?@              8@      �?      @              @      �?      @      �?                      @      <@      3@      "@      *@       @      �?      @              @      �?       @      �?       @                      �?       @              �?      (@              &@      �?      �?      �?                      �?      3@      @      3@       @      .@              @       @      @              �?       @      �?                       @              @     �n@      J@      l@      C@     �b@      *@     �C@              \@      *@      4@      @              @      4@      @      0@              @      @      @              �?      @              @      �?              W@      @      @       @      @              �?       @               @      �?              V@      @      U@       @      Q@              0@       @              �?      0@      �?      .@              �?      �?              �?      �?              @       @               @      @             @R@      9@     @R@      4@      @             �P@      4@      N@      .@      &@      @      &@      @       @      @      �?              �?      @              @      �?              "@                       @     �H@       @     �C@       @      .@              8@       @              �?      8@      �?      5@              @      �?              �?      @              $@      @      @      @      @      @      @      �?       @              �?      �?      �?                      �?               @              @      @              @      @      @              @      @      @      @      @      �?       @      �?       @                      �?      �?                       @               @              @      5@      ,@              @      5@      &@      5@      "@      1@      "@      �?      @      �?                      @      0@      @      .@      �?      ,@              �?      �?              �?      �?              �?      @              @      �?              @                       @      Q@     �q@      <@      C@      <@      >@      @              9@      >@      3@      >@      (@      @      @      @      @       @      @              �?       @              �?      �?      �?      �?                      �?              @      @              @      8@      @      6@      @      ,@      @      $@      @              �?      $@              @      �?      @              @      �?       @      �?                       @              @               @      @       @      @                       @      @                       @      D@     �n@      3@      l@      (@      M@      "@     �L@       @     �D@       @      ;@              (@       @      .@      �?              �?      .@      �?      @      �?       @               @      �?                      �?              (@              ,@      @      0@      �?      ,@      �?      @              @      �?                       @      @       @      @                       @      @      �?       @              �?      �?              �?      �?              @     �d@      @     �d@      @     �U@      @     @S@       @      S@       @      ;@      �?      9@      �?      "@              @      �?      @      �?                      @              0@      �?       @      �?                       @             �H@      �?      �?              �?      �?              @      $@       @      �?              �?       @              �?      "@              "@      �?                     �S@      �?       @      �?                       @      5@      5@      1@      5@      *@      $@      *@      @      *@      �?      &@               @      �?              �?       @                      @              @      @      &@       @      &@              @       @      @       @      �?       @                      �?              @       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK݅�h}�BX0         ~                    �?�#i����?�           ��@       3                    �?<=�h)W�?           �{@       $       	          ����?�r*e���?\            �b@       	                   @E@��C����?:            �W@                            E@���N8�?             5@                           @D@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     1@
       #                    �?rr�J��?+            �R@                          @Z@�m����?#            �M@������������������������       �                     @                          `_@��k��?             �J@������������������������       �                     &@                           @F@և���X�?             E@                          @b@ףp=
�?             $@                           a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           d@     ��?             @@                           �?r�q��?             8@������������������������       �                     @                          �_@������?
             1@              	            �?X�<ݚ�?             "@                          �^@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @       "                   `a@      �?              @        !                    �J@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@%       *                   Pl@f1r��g�?"            �J@&       '                    @Q@�FVQ&�?            �@@������������������������       �                     >@(       )                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?+       ,                   �^@�z�G��?             4@������������������������       �                      @-       .                   �n@�<ݚ�?             2@������������������������       �                     @/       0                   xu@��S�ۿ?	             .@������������������������       �                     &@1       2       	             �?      �?             @������������������������       �                     �?������������������������       �                     @4       ;                    @F@���@��?�            �r@5       :       	             @�x�E~�?5            @V@6       9                   �a@�|���?4             V@7       8                    @B@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �        -            @S@������������������������       �                     �?<       k       	          pff�?P;8����?�            �i@=       `                    �?p`q�q��?e            �c@>       E                    �?     ��?S             `@?       D                    _@���.�6�?$             G@@       C                     L@     ��?             0@A       B                   �V@�r����?             .@������������������������       �                      @������������������������       �        
             *@������������������������       �                     �?������������������������       �                     >@F       _                     P@��P���?/            �T@G       ^                   ht@P�~D&�?'            �P@H       K                   @[@     ��?&             P@I       J                    @I@և���X�?             @������������������������       �                     @������������������������       �                     @L       S                   pa@F�t�K��?#            �L@M       N                    @�>����?             ;@������������������������       �                     5@O       R                   �r@�q�q�?             @P       Q                    ^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @T       ]                   Pm@�z�G��?             >@U       \                    �N@�\��N��?             3@V       [                   �b@��.k���?
             1@W       X                    �?��S���?	             .@������������������������       �                     @Y       Z                   �h@�q�q�?             (@������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     &@������������������������       �                     @������������������������       �                     .@a       b                     L@d��0u��?             >@������������������������       �                     "@c       f                   `_@�G��l��?             5@d       e                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @g       j       	          ����?      �?             (@h       i                     N@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @l       m                   �d@`�(c�?            �H@������������������������       �                     (@n       y                   �o@��+��?            �B@o       v       	          ��� @�	j*D�?             :@p       u                    �?��s����?             5@q       t                    �H@�KM�]�?             3@r       s                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             0@������������������������       �                      @w       x                    �O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?z       }                    �?�C��2(�?             &@{       |                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@       �                   �Z@ ]�к��?�             r@�       �                    �?���|���?             &@������������������������       �                     @������������������������       �                     @�       �                    �?^��:��?�            pq@�       �                   �b@rLTAf�?�            �h@�       �                    �?$�{�F"�?s             e@�       �                    �?X�<ݚ�?             2@�       �       	          ����?��S���?             .@�       �                   �r@�<ݚ�?             "@������������������������       �                     @�       �                   �s@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     J@r�q��?             @������������������������       �                     @�       �                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          ����?,I�e���?f            �b@�       �                    @j(���?4            @S@�       �                    �?>A�F<�?3             S@�       �                   �b@f1r��g�?%            �J@�       �                   i@�:�^���?             �F@������������������������       �                     6@�       �                   @_@�㙢�c�?             7@�       �       	          ����?�����H�?             2@�       �                    @K@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@�       �                   0n@���Q��?             @�       �                   @`@�q�q�?             @�       �                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     @�       �                   @^@��+7��?             7@�       �                    �N@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �]@�t����?
             1@������������������������       �                     @�       �                   a@z�G�z�?             $@�       �                   P`@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   @^@�?�|�?2            �R@�       �       	          ��� @�KM�]�?             3@�       �                    �L@����X�?             @������������������������       �                     @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@������������������������       �        '            �K@�       �       	          033�?�q�q�?             >@�       �                    �?�S����?             3@�       �                    h@���!pc�?             &@������������������������       �                     �?�       �                   pn@z�G�z�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �\@���|���?             &@������������������������       �                      @�       �                   �q@X�<ݚ�?             "@�       �                   �c@և���X�?             @�       �                    @B@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?P���Q�?0             T@������������������������       �        (            �P@�       �                   �`@����X�?             ,@�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @�       �       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       `u@     �x@     �q@     �c@      K@     �W@      G@     �H@      �?      4@      �?      @              @      �?                      1@     �F@      =@      >@      =@      @              8@      =@              &@      8@      2@      �?      "@      �?       @               @      �?                      @      7@      "@      4@      @      @              *@      @      @      @      @      @      @                      @              �?       @              @      @      @      �?      @                      �?              @      .@               @     �F@       @      ?@              >@       @      �?       @                      �?      @      ,@       @              @      ,@      @              �?      ,@              &@      �?      @      �?                      @      m@      P@     �U@       @     �U@      �?      $@      �?              �?      $@             @S@                      �?      b@      O@     �_@      @@     �Z@      5@     �E@      @      *@      @      *@       @               @      *@                      �?      >@              P@      2@     �H@      2@     �H@      .@      @      @              @      @              G@      &@      9@       @      5@              @       @      �?       @      �?                       @      @              5@      "@      $@      "@       @      "@       @      @      @              @      @      @                      @               @       @              &@                      @      .@              3@      &@      "@              $@      &@      �?       @      �?                       @      "@      @      �?      @      �?                      @       @              3@      >@              (@      3@      2@      2@       @      1@      @      1@       @      �?       @               @      �?              0@                       @      �?      @              @      �?              �?      $@      �?      �?      �?                      �?              "@      L@     @m@      @      @              @      @             �H@     �l@     �F@     @c@      9@      b@       @      $@       @      @      @       @      @              �?       @               @      �?              �?      @              @      �?       @               @      �?                      @      1@     �`@      .@      O@      ,@      O@       @     �F@      @     �D@              6@      @      3@       @      0@       @      @              @       @                      &@       @      @       @      �?      �?      �?              �?      �?              �?                       @      @      @      @                      @      @      1@      @       @      @                       @       @      .@              @       @       @       @      @       @                      @              @      �?               @      R@       @      1@       @      @              @       @      �?       @                      �?              (@             �K@      4@      $@      0@      @       @      @              �?       @       @      @              @       @              �?      @      �?      @                      �?       @              @      @               @      @      @      @      @      @      �?              �?      @                       @               @      @      S@             �P@      @      $@      @      @              @      @              �?      @      �?      @      �?                      @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK텔h}�B�3         l                   �`@�/�$�y�?�           ��@       E                    �?R�����?�            @v@              	          ����?H%u��?�            @o@                           @O@(���@��?             �G@                           �?�n_Y�K�?            �C@������������������������       �                     @                          �e@">�֕�?            �A@       	                    �?@�0�!��?
             1@������������������������       �                     *@
                           [@      �?             @������������������������       �                     �?������������������������       �                     @                          �h@X�<ݚ�?             2@������������������������       �                     @                           �?�q�q�?             .@                          �p@z�G�z�?             $@                           �?      �?              @                          @Z@      �?             @                           �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           `@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @       <                   8s@��ؠ���?�            `i@        7                   P`@�;Y�&��?q            @f@!       (                    �?���U�?j            `e@"       #                   @]@�<ݚ�?	             "@������������������������       �                     @$       %                    `@�q�q�?             @������������������������       �                     @&       '       	          433�?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       0       	          033@F|/ߨ�?a            @d@*       /                    �L@@x�5?�?W             b@+       ,                    @L@�k~X��?,             R@������������������������       �        &             P@-       .                   �^@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �        +             R@1       6                   �\@r�q��?
             2@2       3                    �?�q�q�?             "@������������������������       �                     @4       5                     M@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     "@8       ;                   0i@և���X�?             @9       :       	             @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @=       @       	             �?�+e�X�?             9@>       ?                   ��@z�G�z�?             @������������������������       �                     @������������������������       �                     �?A       B                    �?ףp=
�?             4@������������������������       �                     ,@C       D                    @Q@�q�q�?             @������������������������       �                     @������������������������       �                      @F       Q                    �?      �?>            �Z@G       P                    �?b�h�d.�?            �A@H       M                   v@<���D�?            �@@I       L                   �p@ 	��p�?             =@J       K                   �n@�r����?	             .@������������������������       �                     *@������������������������       �                      @������������������������       �                     ,@N       O                   �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @R       c                    �?��U��?+            �Q@S       b                    @      �?             C@T       _       	             �?4���C�?            �@@U       X                   @_@�q�q�?             8@V       W                   `X@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @Y       Z                    �?�r����?             .@������������������������       �                     @[       ^       	          ����?      �?              @\       ]                    �N@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @`       a                    �P@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @d       e                   @\@6YE�t�?            �@@������������������������       �                      @f       k                   P`@��a�n`�?             ?@g       j                     N@���!pc�?             &@h       i                   �_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     4@m       �                    �?������?�            �w@n       �       	          ����?�7����?\            �a@o       p                   @E@�^�����?*             O@������������������������       �                     @q       �                   (q@\�����?%            �K@r       w                    i@">�֕�?            �A@s       v                   @_@��
ц��?             *@t       u                    b@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @x       y                    �?"pc�
�?             6@������������������������       �                      @z                           �?����X�?             ,@{       ~                   pf@�	j*D�?
             *@|       }                    �I@      �?	             (@������������������������       �                     "@������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �_@      �?             4@������������������������       �                     &@�       �                   �d@X�<ݚ�?             "@�       �                    s@�q�q�?             @������������������������       �                     �?�       �                   �s@z�G�z�?             @������������������������       �                     @�       �                     K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �G@�+ت�M�?2            �S@�       �                    @F@���|���?	             &@�       �                   e@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   �c@l��\��?)             Q@�       �                    �?h㱪��?            �K@�       �       	          `ff�?      �?             0@������������������������       �                     (@�       �                   �a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                    �C@�       �       	          ����?�	j*D�?
             *@�       �                    @J@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?�����H�?             "@������������������������       �                     @�       �                    �L@z�G�z�?             @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�P�����?�            �m@�       �                   @g@ ,��-�?H            �]@�       �                   p@؞�z�̼?G            @]@������������������������       �        -            @S@�       �                    �?z�G�z�?             D@�       �                     C@������?            �B@�       �                    �A@���Q��?             @�       �                   @`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    @L@      �?             @@������������������������       �                     =@�       �                    q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �c@^;|��?M            �]@�       �                    �?�z�G��?             $@�       �                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `c@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �k@:��Z��?F            @[@�       �                    �L@��E�B��?            �G@�       �       	          033�?��p\�?            �D@�       �                   �c@������?             B@�       �                   Pc@��S�ۿ?             .@������������������������       �        
             ,@������������������������       �                     �?������������������������       �        	             5@�       �                    i@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                   Pm@¦	^_�?,             O@�       �       	          033@      �?
             ,@�       �                    _@�z�G��?             $@������������������������       �                     @�       �       	          ����?և���X�?             @�       �                   �l@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�q�q��?"             H@�       �                   `a@8�Z$���?            �C@�       �       	             �?h�����?             <@������������������������       �                     7@�       �       	          ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    d@�eP*L��?	             &@�       �                   �d@���Q��?             $@�       �                   �o@�q�q�?             @������������������������       �                     �?�       �                   �r@z�G�z�?             @������������������������       �                     @�       �                   t@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �G@X�<ݚ�?             "@������������������������       �                     @�       �       	          033�?�q�q�?             @������������������������       �                     @������������������������       �                      @�t�b�$     h�h(h+K ��h-��R�(KK�KK��h^�B�        t@     �y@     �T@     q@      >@     �k@      .@      @@      .@      8@      @              &@      8@      @      ,@              *@      @      �?              �?      @               @      $@      @              @      $@       @       @      �?      @      �?      @      �?      �?              �?      �?                       @              @      �?      �?              �?      �?              @       @      @                       @               @      .@     �g@      "@      e@      @     �d@       @      @              @       @      @              @       @      �?              �?       @              @     �c@      �?     �a@      �?     �Q@              P@      �?      @              @      �?                      R@      @      .@      @      @              @      @      @      @                      @              "@      @      @      @      �?      @                      �?              @      @      3@      @      �?      @                      �?       @      2@              ,@       @      @              @       @             �J@     �J@      =@      @      =@      @      ;@       @      *@       @      *@                       @      ,@               @       @               @       @                       @      8@     �G@      3@      3@      3@      ,@      1@      @      @      @              @      @              *@       @      @              @       @      @       @      @                       @       @               @      @              @       @                      @      @      <@       @              @      <@      @       @      @      �?              �?      @                      @              4@     �m@     �a@     �C@     �Y@      =@     �@@              @      =@      :@      8@      &@      @      @       @      @       @                      @      @              2@      @       @              $@      @      "@      @      "@      @      "@                      @              �?      �?              @      .@              &@      @      @       @      @      �?              �?      @              @      �?      �?              �?      �?              @              $@     @Q@      @      @       @      @              @       @               @              @      O@       @     �J@       @      ,@              (@       @       @       @                       @             �C@      @      "@      @      �?              �?      @              �?       @              @      �?      @      �?      �?      �?                      �?              @     �h@     �C@     �[@       @     �[@      @     @S@             �@@      @     �@@      @       @      @       @       @               @       @                      �?      ?@      �?      =@               @      �?              �?       @                      @              �?      V@      ?@      @      @      �?      @              @      �?               @      @              @       @             @U@      8@     �D@      @      C@      @     �A@      �?      ,@      �?      ,@                      �?      5@              @       @               @      @              @      @              @      @              F@      2@      @      @      @      @      @              @      @      �?      @      �?                      @      @                      @     �B@      &@     �@@      @      ;@      �?      7@              @      �?              �?      @              @      @      @      @       @      @      �?              �?      @              @      �?      �?      �?                      �?      @                      �?      @      @              @      @       @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KKۅ�h}�B�/         V                   �`@���
%�?�           ��@       3                    �?�ڳ�$��?�            �t@       2                   pz@$]^z���?�             m@       1                    �R@�����?�            �l@                           �?�W�a=�?�            �l@              	          ����?�GN�z�?(            �P@       
                    �?���3�E�?             J@       	                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @                           �?�5��
J�?             G@              	          ����?�S����?             C@              	          ���ܿz�G�z�?             >@������������������������       �                     �?                           [@V�a�� �?             =@                          �_@�q�q�?             "@                          �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �V@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             4@������������������������       �                      @                           �L@      �?              @������������������������       �                      @                          �`@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@       .                   xt@Ћ����?k            �d@        '                   �b@�{���l�?f            �c@!       &       	          ����? ����?R            @`@"       #       	          833�? 	��p�?             =@������������������������       �                     5@$       %                   `^@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �        C            @Y@(       -       	             �?�>����?             ;@)       *                    �?���Q��?             @������������������������       �                      @+       ,                   �[@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     6@/       0                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?4       9                    �?     ��?>             X@5       8                   �Z@��S�ۿ?             .@6       7                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             *@:       U                    �?:~=�P�?2            @T@;       T                    `@�U���?&             O@<       I                    �?���dQ'�?#            �L@=       B                    �?�q�q�?             2@>       ?                     Q@z�G�z�?             @������������������������       �                     @@       A                     R@      �?              @������������������������       �                     �?������������������������       �                     �?C       H                    @K@8�Z$���?
             *@D       E                   `X@�q�q�?             @������������������������       �                     �?F       G                   �S@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @J       S                    @x�����?            �C@K       L                   �m@�MI8d�?            �B@������������������������       �                     7@M       N                   �U@և���X�?             ,@������������������������       �                     @O       R                   �`@���!pc�?             &@P       Q                   @_@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     3@W       f                   �O@>n�T��?�            `y@X       a                    �?؇���X�?             <@Y       `                    �?�C��2(�?             6@Z       [                     H@      �?              @������������������������       �                     @\       ]                    �?���Q��?             @������������������������       �                      @^       _       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             ,@b       c                   �b@�q�q�?             @������������������������       �                      @d       e                    `@      �?             @������������������������       �                      @������������������������       �                      @g       �       	          pff�?�I�E��?�            �w@h       �                    @L@�X3����?�            `p@i       �                    �?������?�             j@j       �                    @I@�!�I�*�?x            �g@k       �                   �p@�}�x�m�?O            �^@l       �                    �?��l��??            @X@m       n                   `b@��a�n`�?<            @W@������������������������       �                     4@o       �                    �?0�й���?1            @R@p       w                    @G@��ɉ�?*            @P@q       v                    �?�IєX�?             �I@r       u                    �?���Q��?             @s       t                   �f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     G@x       y                   @c@և���X�?
             ,@������������������������       �                     @z       {                     H@���!pc�?             &@������������������������       �                     �?|                          �p@�z�G��?             $@}       ~                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?      �?             @�       �                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?$��m��?             :@�       �                   �r@�n_Y�K�?             *@������������������������       �                      @������������������������       �                     @�       �                    �?$�q-�?
             *@������������������������       �        	             (@������������������������       �                     �?�       �                    �?�\=lf�?)            �P@�       �                    f@ qP��B�?            �E@������������������������       �                     E@������������������������       �                     �?������������������������       �                     8@�       �                   �^@D�n�3�?             3@�       �                    c@      �?              @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?"pc�
�?             &@������������������������       �                      @������������������������       �                     "@�       �                   �d@Fmq��?%            �J@�       �                   �e@��H�}�?#             I@������������������������       �                     @�       �       	          pff�?�û��|�?              G@�       �                   �_@�c�Α�?             =@�       �                   @n@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?"pc�
�?             6@������������������������       �                     @�       �                    �?������?             .@�       �                   `a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �r@r�q��?             (@�       �                    �?�C��2(�?
             &@������������������������       �                     "@�       �                   �h@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   Pd@j���� �?
             1@�       �                    @N@�θ�?             *@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   pc@�c�Α�?@             ]@�       �                    �?&^�)b�?-            �U@�       �                    �?և���X�?             5@�       �                     K@"pc�
�?             &@�       �                   Pn@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                   �Z@����?"            @P@������������������������       �                     �?�       �       	          ����?     �?!             P@�       �                    j@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0c@�]0��<�?            �N@�       �                   `a@ _�@�Y�?             M@�       �                     P@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     H@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	             @��S���?             >@�       �                   �`@���!pc�?             6@�       �                    �L@؇���X�?	             ,@������������������������       �                     "@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       0s@     �z@      O@     �p@      7@      j@      6@      j@      5@      j@      .@     �I@      .@     �B@      @       @      @                       @      &@     �A@      @      @@      @      8@              �?      @      7@      @      @      �?       @               @      �?              @      �?              �?      @                      4@               @      @      @               @      @      �?      @                      �?              ,@      @     �c@      @      c@       @      `@       @      ;@              5@       @      @              @       @                     @Y@       @      9@       @      @               @       @      �?              �?       @                      6@       @      @       @                      @      �?              �?             �C@     �L@      ,@      �?      �?      �?              �?      �?              *@              9@      L@      9@     �B@      4@     �B@      (@      @      �?      @              @      �?      �?      �?                      �?      &@       @      @       @              �?      @      �?              �?      @              @               @      ?@      @      ?@              7@      @       @      @              @       @      @       @               @      @                      @       @              @                      3@     �n@      d@      @      8@       @      4@       @      @              @       @      @               @       @      �?              �?       @                      ,@       @      @               @       @       @               @       @              n@      a@      j@     �J@      f@      @@      e@      5@     �Y@      4@     �U@      &@      U@      "@      4@              P@      "@      L@      "@      H@      @       @      @       @      �?              �?       @                       @      G@               @      @              @       @      @      �?              @      @      @      @      @                      @      @               @               @       @      �?       @               @      �?              �?              1@      "@      @       @               @      @              (@      �?      (@                      �?     �P@      �?      E@      �?      E@                      �?      8@               @      &@      @       @      �?       @               @      �?              @               @      "@       @                      "@      @@      5@      @@      2@      @              <@      2@      5@       @      @      @      @                      @      2@      @      @              &@      @      �?       @      �?                       @      $@       @      $@      �?      "@              �?      �?      �?                      �?              �?      @      $@      @      $@              @      @      @              @      @              @                      @      @@      U@      0@     �Q@      (@      "@       @      "@       @       @       @                       @              @      $@              @     �N@      �?              @     �N@      �?       @      �?                       @       @     �M@      �?     �L@      �?      "@              "@      �?                      H@      �?       @      �?                       @      0@      ,@      0@      @      (@       @      "@              @       @      @                       @      @      @              @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK녔h}�Bh3         �       	          033�?�r,��?�           ��@       m                    �?H;N	�	�?�             x@                          @E@`Y�K�?�            �s@       	                    �?^������?            �A@              	          ����?�LQ�1	�?             7@������������������������       �        
             2@              	          833�?���Q��?             @������������������������       �                     @������������������������       �                      @
                           ^@      �?             (@������������������������       �                      @                           @I@      �?             @������������������������       �                      @              	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?       >                    �?�����?�            Pq@       3                   8q@�D����?0             U@       .                   �a@
��[��?&            @P@       %                   �b@^l��[B�?!             M@                          �j@؇���X�?             E@                          �`@���7�?             6@                           �?$�q-�?             *@                           `@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                      @������������������������       �                     "@                           k@      �?             4@������������������������       �                      @                            �?r�q��?             2@������������������������       �                      @!       "                    �?      �?
             0@������������������������       �                     ,@#       $                    l@      �?              @������������������������       �                     �?������������������������       �                     �?&       '                   �c@     ��?
             0@������������������������       �                     @(       -       	             �?      �?             (@)       ,                   `i@�q�q�?             "@*       +                   �f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @/       0                   �`@����X�?             @������������������������       �                      @1       2                    �?���Q��?             @������������������������       �                     @������������������������       �                      @4       9                   Hw@�S����?
             3@5       6                    �F@��S�ۿ?             .@������������������������       �                     @7       8                    a@      �?              @������������������������       �                     �?������������������������       �                     @:       ;                     C@      �?             @������������������������       �                     �?<       =                   8|@�q�q�?             @������������������������       �                      @������������������������       �                     �??       X                    @L@����ڽ?�             h@@       O                   �q@(;L]n�?e            �b@A       B                   �`@     ��?W             `@������������������������       �        B            �X@C       D                    �? 	��p�?             =@������������������������       �        
             1@E       F                   �`@r�q��?             (@������������������������       �                     �?G       H                    �G@�C��2(�?
             &@������������������������       �                     @I       J                   0d@r�q��?             @������������������������       �                     @K       L                   @a@�q�q�?             @������������������������       �                     �?M       N                    �?      �?              @������������������������       �                     �?������������������������       �                     �?P       W                    @��2(&�?             6@Q       V                    �?P���Q�?             4@R       U                    �?      �?             @S       T                    d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             0@������������������������       �                      @Y       Z                    �?�T|n�q�?            �E@������������������������       �                     $@[       h                    �?�'�`d�?            �@@\       ]                    �L@\-��p�?             =@������������������������       �                     �?^       c                    �M@ �Cc}�?             <@_       b       	          ����?z�G�z�?             $@`       a                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?d       e                   ht@�X�<ݺ?             2@������������������������       �        
             0@f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?i       l                   Pa@      �?             @j       k                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @n       �                    �?^H���+�?.            �R@o       ~                   �b@x��}�?!            �K@p       u                   pb@�:�^���?            �F@q       r                   �p@      �?             @@������������������������       �                     >@s       t                    �?      �?              @������������������������       �                     �?������������������������       �                     �?v       w                    �?�θ�?             *@������������������������       �                     �?x       }                   �c@      �?             (@y       |                   �b@���Q��?             @z       {                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @       �                   @j@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    ]@�����?             3@������������������������       �                     @�       �                    �?��
ц��?
             *@�       �                    �?���|���?             &@�       �                   �b@�<ݚ�?             "@�       �                   Xp@      �?              @�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?д>��C�?�            �u@�       �                   �[@���B��?@            @Y@������������������������       �                     &@�       �                   �]@b�2�tk�?8            �V@�       �                    �D@�����H�?             "@�       �                     C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �L@�q�q�?2            @T@�       �                    m@��
ц��?            �C@�       �                   �b@$��m��?             :@�       �       	             �?$�q-�?
             *@������������������������       �                     �?������������������������       �        	             (@�       �                    U@�n_Y�K�?             *@������������������������       �                      @�       �       	          ����?���!pc�?             &@������������������������       �                     @������������������������       �                      @�       �                   (p@$�q-�?
             *@������������������������       �                      @�       �       	          ���@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?؇���X�?             E@�       �                    @V�a�� �?             =@�       �                   @[@PN��T'�?             ;@������������������������       �                     @�       �                   `v@ �q�q�?             8@������������������������       �                     6@�       �       	          ���@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@�       �                    @G@`Pp�I�?�            �n@�       �                    �?�c�Α�?             =@�       �                    @C@      �?             <@������������������������       �                     "@�       �                   �m@p�ݯ��?             3@�       �                   �`@��
ц��?	             *@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �?���qh�?�            @k@�       �                   `c@�θ�?             :@�       �                    a@���Q��?
             .@�       �                   @[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       	          033�?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     &@�       �                    @p�q��?{             h@�       �                    V@���g�?z            �g@������������������������       �                     �?�       �                   P`@�# ��?y            �g@�       �                   �`@\#r��?+            �N@�       �                    �?��E�B��?!            �G@�       �                    �?�n`���?             ?@�       �       	          033@؇���X�?             <@�       �                    �?H%u��?             9@������������������������       �                     "@�       �                    @L@     ��?             0@������������������������       �                     $@�       �                    n@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             0@������������������������       �        
             ,@�       �                    �? qP��B�?N             `@������������������������       �        2            �T@�       �       	          ����?���.�6�?             G@�       �                   �b@R���Q�?             4@������������������������       �        	             *@�       �                   �`@և���X�?             @�       �                     L@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     :@������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h^�B�       �t@     Py@     �p@     @]@     `n@     @Q@      (@      7@      @      4@              2@      @       @      @                       @      "@      @       @              �?      @               @      �?      �?              �?      �?             �l@      G@      I@      A@     �G@      2@     �F@      *@      B@      @      5@      �?      (@      �?      $@      �?              �?      $@               @              "@              .@      @               @      .@      @               @      .@      �?      ,@              �?      �?              �?      �?              "@      @              @      "@      @      @      @      �?      @              @      �?              @              @               @      @               @       @      @              @       @              @      0@      �?      ,@              @      �?      @      �?                      @       @       @              �?       @      �?       @                      �?     �f@      (@      b@      @     �_@       @     �X@              ;@       @      1@              $@       @              �?      $@      �?      @              @      �?      @               @      �?      �?              �?      �?              �?      �?              3@      @      3@      �?      @      �?       @      �?       @                      �?      �?              0@                       @      B@      @      $@              :@      @      9@      @              �?      9@      @       @       @       @      �?       @                      �?              �?      1@      �?      0@              �?      �?      �?                      �?      �?      @      �?      �?      �?                      �?               @      :@      H@      *@      E@      @     �D@      �?      ?@              >@      �?      �?              �?      �?              @      $@              �?      @      "@      @       @      �?       @      �?                       @       @                      @      "@      �?              �?      "@              *@      @      @              @      @      @      @      @       @      @      �?      �?      �?              �?      �?              @                      �?               @               @      N@      r@     �A@     �P@              &@     �A@     �K@       @      �?      �?      �?      �?                      �?      @              ;@      K@      5@      2@      "@      1@      �?      (@      �?                      (@       @      @               @       @      @              @       @              (@      �?       @              @      �?      @                      �?      @      B@      @      7@      @      7@      @              �?      7@              6@      �?      �?      �?                      �?       @                      *@      9@     �k@       @      5@      @      5@              "@      @      (@      @      @              @      @                      @      �?              1@      i@      @      4@      @      "@      @      �?              �?      @               @       @               @       @                      &@      &@     �f@      $@     �f@      �?              "@     �f@      @     �K@      @     �D@      @      9@      @      8@      @      6@              "@      @      *@              $@      @      @      @                      @      �?       @               @      �?               @      �?              �?       @                      0@              ,@      @     �_@             �T@      @     �E@      @      1@              *@      @      @       @      �?              �?       @              �?      @              @      �?                      :@      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK兔h}�B2         P                   �`@T8���?�           ��@       7       	             �?�f@���?�            �u@                          �a@J!�k���?P             `@                           �? {��e�?!            �J@                          �_@V������?            �B@       	       	             п�KM�]�?             3@                           �N@      �?              @������������������������       �                     �?������������������������       �                     �?
                            E@�IєX�?	             1@������������������������       �                     �?������������������������       �                     0@                           �?      �?             2@                           �?"pc�
�?             &@                          �[@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        
             0@       ,                    �?���=A�?/             S@       +                   (@z�G�z�?"            �K@       *                    �Q@8�Z$���?!             J@                           �?L紂P�?             �I@������������������������       �        	             (@                           �F@:�&���?            �C@������������������������       �                     "@       )                    q@�������?             >@                           �]@�>4և��?             <@                          @Z@���Q��?             @������������������������       �                     @������������������������       �                      @!       "                   �[@�LQ�1	�?             7@������������������������       �                     $@#       &                   �`@�θ�?             *@$       %                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?'       (                    ]@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @-       6                   �s@�q�q�?             5@.       3                   �]@     ��?             0@/       2                   xp@���!pc�?             &@0       1       	          ����?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @4       5                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @8       9                   �Q@�o�s(��?�            �k@������������������������       �                     �?:       E                    �?�2����?�            `k@;       >                    �?���Q��?
             .@<       =                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @?       D       	             @�q�q�?             (@@       C                   �d@z�G�z�?             $@A       B                    �H@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @F       K                   0`@���J��?            �i@G       H                   �c@@~��?q            @f@������������������������       �        \            �b@I       J                     R@h�����?             <@������������������������       �                     ;@������������������������       �                     �?L       M                    �?ȵHPS!�?             :@������������������������       �        	             .@N       O                   �a@���!pc�?             &@������������������������       �                      @������������������������       �                     @Q       �                    �?d��Mܻ�?�            x@R       �                    �?|�{���?]            �`@S       f                    �?X�<ݚ�?J             [@T       e       	          `ff@b�2�tk�?             B@U       V                   `T@     ��?             @@������������������������       �                     @W       b                   �a@>���Rp�?             =@X       _                   �d@      �?             8@Y       Z                    �?�C��2(�?             6@������������������������       �                     $@[       \                   �r@r�q��?             (@������������������������       �                      @]       ^                   c@      �?             @������������������������       �                      @������������������������       �                      @`       a                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?c       d                    c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @g       �                    �?*O���?3             R@h       q                   �b@      �?             C@i       j                   @j@"pc�
�?	             &@������������������������       �                     @k       p       	          tff�?���Q��?             @l       o                   �a@      �?             @m       n       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?r              	          ����?��}*_��?             ;@s       ~                   �r@`�Q��?             9@t       }                   �o@�GN�z�?             6@u       v                   �\@�n_Y�K�?             *@������������������������       �                     @w       |                   l@      �?              @x       {                    a@      �?             @y       z                   Pi@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                      @�       �       	             �?H�V�e��?             A@�       �                   �d@�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                   @M@r�q��?             8@�       �                   �`@�q�q�?             @������������������������       �                     �?�       �                   @Z@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �m@�����?             5@�       �                    �G@r�q��?	             (@�       �                    �D@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                   �[@ 7���B�?             ;@�       �                    ]@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     6@�       �                    @j�q����?�            @o@�       �       	          033�?Vd*�=�?�            �l@�       �                   �a@�����?{            �h@�       �                    �?     ��?             @@�       �                   p@�J�4�?             9@������������������������       �                     .@�       �       	            �?���Q��?             $@�       �                   a@�q�q�?             @������������������������       �                     �?�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    q@      �?             @������������������������       �                      @������������������������       �                      @�       �                   @f@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   h@���*�?h            �d@�       �       	          ����?P%�Ѿ�?f            �d@�       �                   �t@�7�	|��?L             `@������������������������       �        J            �_@�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �Q@b�h�d.�?            �A@������������������������       �                     �?�       �                   �b@��hJ,�?             A@�       �                   �p@      �?             @������������������������       �                      @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �g@��S�ۿ?             >@�       �                    �?�q�q�?             @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   0a@ 7���B�?             ;@������������������������       �                     4@�       �                   m@؇���X�?             @������������������������       �                     @�       �                   xp@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   pn@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?l��[B��?             =@������������������������       �                     @�       �                   �c@�LQ�1	�?             7@�       �                    �?�8��8��?             (@�       �                   �m@�C��2(�?             &@������������������������       �                      @�       �                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    @G@���|���?             &@������������������������       �                     @�       �                    _@և���X�?             @������������������������       �                     �?�       �       	          `ff@�q�q�?             @������������������������       �                     �?�       �                   �d@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   @e@      �?             6@�       �                    �O@b�2�tk�?
             2@�       �                   �[@d}h���?             ,@������������������������       �                      @�       �                   d@�8��8��?             (@������������������������       �                     $@�       �                   pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h^�BP       �t@     @y@      S@     q@      O@     �P@      &@      E@      &@      :@       @      1@      �?      �?              �?      �?              �?      0@      �?                      0@      "@      "@      "@       @      @       @      @                       @      @                      @              0@     �I@      9@      F@      &@      F@       @      F@      @      (@              @@      @      "@              7@      @      7@      @      @       @      @                       @      4@      @      $@              $@      @      �?       @               @      �?              "@      �?              �?      "@                       @              �?              @      @      ,@      @      "@      @       @      @      @              @      @                      @      @      �?      @                      �?              @      ,@     �i@      �?              *@     �i@      "@      @      �?       @      �?                       @       @      @       @       @       @      �?              �?       @                      �?               @      @      i@      �?      f@             �b@      �?      ;@              ;@      �?              @      7@              .@      @       @               @      @             �o@     ``@     �H@     �U@      H@      N@      6@      ,@      6@      $@              @      6@      @      5@      @      4@       @      $@              $@       @       @               @       @               @       @              �?      �?              �?      �?              �?      @              @      �?                      @      :@      G@      3@      3@      "@       @      @              @       @      @      �?      �?      �?              �?      �?               @                      �?      $@      1@       @      1@      @      1@      @       @              @      @      @      �?      @      �?      �?              �?      �?                       @      @                      "@      @               @              @      ;@      @      @              @      @              @      4@       @      �?      �?              �?      �?      �?                      �?       @      3@       @      $@       @      @              @       @                      @              "@      �?      :@      �?      @              @      �?                      6@     �i@     �F@     @h@      A@     �f@      3@      6@      $@      5@      @      .@              @      @      @       @      �?              @       @               @      @               @       @               @       @              �?      @      �?                      @     �c@      "@     �c@      @      `@      �?     �_@              �?      �?              �?      �?              =@      @              �?      =@      @      �?      @               @      �?      �?      �?                      �?      <@       @       @      �?      �?      �?              �?      �?              �?              :@      �?      4@              @      �?      @               @      �?              �?       @              �?       @      �?                       @      ,@      .@      @               @      .@      �?      &@      �?      $@               @      �?       @      �?                       @              �?      @      @      @              @      @      �?               @      @              �?       @      @       @                      @      &@      &@      @      &@      @      &@       @              �?      &@              $@      �?      �?              �?      �?              @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        hDK
hEKhFh(h+K ��h-��R�(KK��h^�C              �?�t�bhRhchMC       ���R�hgKhhhkK
h(h+K ��h-��R�(KK��hM�C       �t�bK��R�}�(hKhuK�hvh(h+K ��h-��R�(KK煔h}�B�2         �                    �?�[��N�?�           ��@       e       	          ����? XөM"�?           �y@       2                    �?�t%Q��?�            �r@                           �A@fK!���?:            �V@������������������������       �                     @                          `_@      �?8             V@                           �?�㙢�c�?             7@       	                     E@������?             1@������������������������       �                      @
                          �h@�r����?
             .@                          �_@$�q-�?             *@������������������������       �                     @                           �J@r�q��?             @������������������������       �                     �?������������������������       �                     @                           @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       #                   �b@�n_Y�K�?'            @P@              	          �����@�0�!��?             A@������������������������       �                      @                           �?      �?             @@������������������������       �                     @                             O@PN��T'�?             ;@              	          ����?�8��8��?
             8@                          �j@؇���X�?             ,@������������������������       �                     "@                          �^@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@!       "                   n@�q�q�?             @������������������������       �                     �?������������������������       �                      @$       )                   �c@���@M^�?             ?@%       &                    �?�����H�?             "@������������������������       �                     @'       (                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @*       +                   `i@      �?             6@������������������������       �                     @,       -                   q@ҳ�wY;�?             1@������������������������       �                      @.       /                    �D@�q�q�?             "@������������������������       �                     @0       1                    �?      �?             @������������������������       �                     @������������������������       �                     @3       d                   �g@T�fU���?{             j@4       Y                    @ ���g=�?z            �i@5       L                    @L@dP-���?p            �g@6       =                    �?x�Y��?\            `c@7       8                   �o@�(\����?2             T@������������������������       �        $            �M@9       <                   �a@�����?             5@:       ;                   �[@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     1@>       ?                    �?��S�ۿ?*            �R@������������������������       �                     &@@       A                    @G@     p�?#             P@������������������������       �                     >@B       C                   @[@��hJ,�?             A@������������������������       �                     @D       K       	          ����?`Jj��?             ?@E       F                   pm@(;L]n�?             >@������������������������       �        
             3@G       H                    �?�C��2(�?             &@������������������������       �                      @I       J                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?M       T                    �?���!pc�?            �@@N       O                    �L@�+e�X�?             9@������������������������       �                     @P       S                   �c@��2(&�?             6@Q       R                   ht@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                      @U       X                   `c@      �?              @V       W                    @P@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?Z       c                    �?D�n�3�?
             3@[       \                    �?��S���?             .@������������������������       �                     @]       b                   �c@�q�q�?             (@^       a                    �?�����H�?             "@_       `       	          @33�?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @f       �                   �r@������?M            �[@g       r                    �?r֛w���?B            @W@h       q                    �?      �?             H@i       j                   d@�LQ�1	�?             7@������������������������       �                      @k       p                    @K@���N8�?             5@l       m                   �`@r�q��?             @������������������������       �                     @n       o       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             .@������������������������       �                     9@s       t                    [@��S���?#            �F@������������������������       �                     @u       z                    �?�p ��?             �D@v       w                   0c@�C��2(�?	             &@������������������������       �                     @x       y                    �H@z�G�z�?             @������������������������       �                     �?������������������������       �                     @{       �       	             @d��0u��?             >@|       �                   �o@�\��N��?             3@}       �       	          033�?X�Cc�?             ,@~       �                     L@z�G�z�?             @       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	          ����?�����H�?             "@������������������������       �                     @�       �                   `g@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   @L@�C��2(�?             &@�       �       	          `ff@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                     Q@�����H�?             2@�       �                    �D@�IєX�?
             1@�       �                   �v@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@������������������������       �                     �?�       �                    �?��k�D�?�            0t@�       �                   @d@X����?�            `o@�       �                    �?,��w�?�            �n@�       �                    f@��8���?t             h@�       �                   `[@���8��?q            `g@�       �                   ``@���J��?            �I@�       �                    @L@���N8�?             5@������������������������       �                     1@�       �                    �L@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     >@�       �       	          ����?ДX��?T             a@�       �       	          033�?��|��?.            �S@�       �                   �[@4և����?#             L@�       �                   @_@      �?             @������������������������       �                     �?�       �                   xp@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?0G���ջ?              J@�       �                   pb@��Y��]�?            �D@������������������������       �                     A@�       �                    @I@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?"pc�
�?             &@������������������������       �                     �?�       �                   �l@ףp=
�?             $@������������������������       �                     @�       �                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @_@���!pc�?             6@������������������������       �                     &@�       �                    �?�eP*L��?             &@�       �                   �i@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�8���?&             M@�       �                    �M@��<b�ƥ?             G@������������������������       �                     <@�       �                   �Y@�X�<ݺ?	             2@������������������������       �                     �?������������������������       �                     1@�       �                   �_@r�q��?	             (@������������������������       �                      @������������������������       �                     $@�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        '             K@�       �                    �?���Q��?             @�       �                     K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?*O���?&             R@�       �       	          033�?��B����?             J@�       �                    �L@����X�?            �A@�       �                    I@�IєX�?	             1@������������������������       �                     �?������������������������       �                     0@�       �                    �N@      �?
             2@�       �                   �d@�n_Y�K�?             *@�       �       	          @33�?z�G�z�?             $@�       �                   ``@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          433�?z�G�z�?             @�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             1@�       �                   �`@P���Q�?
             4@������������������������       �        	             3@������������������������       �                     �?�t�b��      h�h(h+K ��h-��R�(KK�KK��h^�Bp       �s@     Pz@     �p@      b@     `l@     @R@      F@     �G@              @      F@      F@      @      3@      @      *@       @               @      *@      �?      (@              @      �?      @      �?                      @      �?      �?      �?                      �?              @      D@      9@      <@      @               @      <@      @      @              7@      @      6@       @      (@       @      "@              @       @      @                       @      $@              �?       @      �?                       @      (@      3@      �?       @              @      �?       @      �?                       @      &@      &@              @      &@      @       @              @      @              @      @      @              @      @             �f@      :@     �f@      8@     �e@      0@     �b@      @     �S@       @     �M@              3@       @       @       @               @       @              1@             �Q@      @      &@             �M@      @      >@              =@      @              @      =@       @      =@      �?      3@              $@      �?       @               @      �?              �?       @                      �?      8@      "@      3@      @              @      3@      @      3@      �?      3@                      �?               @      @      @      @       @      @                       @              �?      &@       @      @       @      @              @       @      �?       @      �?      @              @      �?                      @      @              @                       @      D@     �Q@      8@     @Q@      @     �F@      @      4@       @              �?      4@      �?      @              @      �?      �?      �?                      �?              .@              9@      5@      8@              @      5@      4@      $@      �?      @              @      �?              �?      @              &@      3@      $@      "@      "@      @      �?      @      �?      �?              �?      �?                      @       @      �?      @              @      �?              �?      @              �?      @              @      �?              �?      $@      �?       @               @      �?                       @      0@       @      0@      �?      �?      �?      �?                      �?      .@                      �?      G@     Pq@      4@     �l@      1@     �l@      1@     �e@      .@     �e@      �?      I@      �?      4@              1@      �?      @      �?                      @              >@      ,@     �^@      &@     �P@      @     �I@       @       @      �?              �?       @      �?                       @      @     �H@      �?      D@              A@      �?      @      �?                      @       @      "@      �?              �?      "@              @      �?       @      �?                       @      @      0@              &@      @      @      @      @      @                      @      @              @     �K@      �?     �F@              <@      �?      1@      �?                      1@       @      $@       @                      $@       @      @              @       @                      K@      @       @      @      �?              �?      @                      �?      :@      G@      9@      ;@      9@      $@      0@      �?              �?      0@              "@      "@       @      @       @       @      @       @               @      @              @                      @      �?      @      �?      �?              �?      �?                      @              1@      �?      3@              3@      �?        �t�bubhhubehhub.